library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package data16_pkg is

	type ram_type is array (0 to 2*140-1) of std_logic_vector(15 downto 0);
	constant data16 : ram_type :=(
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"eada",	x"0000",	
												x"d125",	x"0000",	x"0000",	x"0000",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"0004",	x"000a",	
												x"c313",	x"1cc4",	x"4944",	x"6250"
										);
end data16_pkg;