library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package data32_pkg is

	type ram_type is array (0 to 18479) of std_logic_vector(31 downto 0);
	constant data32 : ram_type :=(
					x"00be11e2",	x"0000008c",	x"20111213",	x"0000eada",	
					x"0000d125",	x"00000000",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"000a0004",	x"1cc4c313",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0001002e",	x"06d006a5",	x"069f06a5",	
					x"068c06a4",	x"06a4069e",	x"069406ae",	x"068b06af",	
					x"06d40705",	x"06cf06ad",	x"06d306d1",	x"06f206d9",	
					x"06e606f8",	x"06eb06b4",	x"06c806e6",	x"070c0703",	
					x"070806f2",	x"06f606b3",	x"06c206c3",	x"06e206ee",	
					x"070206d9",	x"06d906e5",	x"06d406c2",	x"06de06f8",	
					x"06fc06e1",	x"06e506a2",	x"06c706e1",	x"06d806de",	
					x"06d306f1",	x"06f6071f",	x"06c906bc",	x"06e106f3",	
					x"06cd0706",	x"06e4067b",	x"0001102e",	x"069e0685",	
					x"069f06b1",	x"06a20667",	x"068d067a",	x"068b06b3",	
					x"06b206b0",	x"06b00696",	x"06b6069c",	x"068d06dd",	
					x"06e806d7",	x"06ce06be",	x"06dd06c5",	x"06cd06ae",	
					x"06bd06cb",	x"06be06c9",	x"06d70678",	x"06c606d7",	
					x"06df06d7",	x"06d606ce",	x"06f406ac",	x"06d206ba",	
					x"06db06dc",	x"06d206bf",	x"06c706b4",	x"06d906fb",	
					x"06e506f8",	x"06eb06fe",	x"070606e9",	x"06f70701",	
					x"07110701",	x"070606ec",	x"06eb06aa",	x"0001202e",	
					x"067e0695",	x"068c0692",	x"069c0676",	x"06800691",	
					x"069606a7",	x"06c106a3",	x"06a306b2",	x"06af069a",	
					x"06c106c5",	x"06d506b6",	x"06d206bf",	x"06d506c0",	
					x"06c306e7",	x"06ef06bc",	x"06b106ac",	x"06ac068e",	
					x"068d06aa",	x"06a106c6",	x"06be06bd",	x"06c306c5",	
					x"06cd06d1",	x"06d806cb",	x"06c806c7",	x"06bc06ae",	
					x"06cd06d1",	x"06cc06d4",	x"06d306e9",	x"06eb06ea",	
					x"06f106ce",	x"06d406c5",	x"069d06dc",	x"06d2065c",	
					x"0001302e",	x"06510668",	x"0672068a",	x"06880694",	
					x"066f0674",	x"065d068c",	x"069b06b0",	x"06a306a0",	
					x"0699067f",	x"067d06c7",	x"06be06c4",	x"06be06ca",	
					x"06c306dc",	x"06b106db",	x"06ad06c5",	x"06c406bf",	
					x"06b70685",	x"069c06be",	x"06c006c3",	x"06c306c1",	
					x"06c606cb",	x"06b506c7",	x"06bb06cf",	x"06bd06d5",	
					x"06bc06bc",	x"06b506ef",	x"06bc06da",	x"06c306f4",	
					x"06db06ec",	x"06cd0705",	x"06cf06f6",	x"06c406f2",	
					x"06cf069d",	x"000a0004",	x"e54900b0",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0002402e",	x"067f06b0",	x"06990693",	
					x"068906a9",	x"069706d9",	x"06a606c5",	x"06ad06ee",	
					x"06d506eb",	x"06cc06ae",	x"06c906eb",	x"06ed06e4",	
					x"06ca06e2",	x"06e506fb",	x"06d606e4",	x"06ee06e8",	
					x"070406f3",	x"06de06ce",	x"06e0070f",	x"071706fc",	
					x"06ed0702",	x"07000710",	x"06f8071b",	x"070a06fe",	
					x"06f906f9",	x"06e806fa",	x"07050713",	x"0706071f",	
					x"07120721",	x"072a072d",	x"06ff073f",	x"071e0733",	
					x"06f6072f",	x"070f06e3",	x"0002502e",	x"06ae06d1",	
					x"06a206d9",	x"06ad06db",	x"06c606ec",	x"06e8070d",	
					x"06f5070e",	x"06f80710",	x"06f70723",	x"0704072c",	
					x"0720073c",	x"0730072a",	x"071b0733",	x"06ea0724",	
					x"072a073f",	x"06ee0731",	x"0702070b",	x"0712072d",	
					x"07130749",	x"0717073d",	x"07230739",	x"071f0740",	
					x"07180745",	x"071d0755",	x"0716073d",	x"0709074a",	
					x"07350770",	x"0739075d",	x"07210774",	x"072d0763",	
					x"0731076f",	x"07260752",	x"070b0700",	x"0002602e",	
					x"06c40715",	x"06dd0713",	x"06d5070a",	x"06fa072d",	
					x"06ea0724",	x"06f60715",	x"06f0072c",	x"06fd072c",	
					x"07080743",	x"07340741",	x"072e073a",	x"073c0768",	
					x"07360757",	x"075f076b",	x"074f076d",	x"073d0743",	
					x"07290774",	x"075b0763",	x"07580773",	x"075a0770",	
					x"0753075d",	x"07530776",	x"0752077f",	x"076f0756",	
					x"07510782",	x"07610781",	x"07420787",	x"0760079a",	
					x"074f07a6",	x"07510782",	x"075a078f",	x"075d0754",	
					x"0002702e",	x"071f075b",	x"071a0731",	x"06e2072d",	
					x"0718077a",	x"07290765",	x"0734078b",	x"075e076d",	
					x"07530752",	x"073b077f",	x"079307ae",	x"078807a6",	
					x"077907b7",	x"075b07a9",	x"07a207c7",	x"077907b3",	
					x"078107ae",	x"078207be",	x"078a07c5",	x"07a307cf",	
					x"078a07ea",	x"07a007d3",	x"07b207c9",	x"079907be",	
					x"07c007bb",	x"07af07ef",	x"07dd0811",	x"07d607fd",	
					x"07e50800",	x"07c10819",	x"07e30821",	x"08020810",	
					x"07ea0630",	x"000a0004",	x"185f43fe",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1003002e",	x"06330644",	x"0661064a",	
					x"0665063b",	x"0651064f",	x"06510693",	x"069a0686",	
					x"066f068e",	x"068e0676",	x"0674066b",	x"06870689",	
					x"0690067c",	x"06a606b2",	x"068e06b1",	x"06cd0692",	
					x"06a3068f",	x"068c0660",	x"0669069d",	x"06a3069b",	
					x"06770681",	x"06920690",	x"069206a9",	x"06a606bc",	
					x"06b50689",	x"06af066c",	x"06a006a6",	x"06a306b8",	
					x"06b506ba",	x"06aa06ad",	x"069606a2",	x"068b06a9",	
					x"068b06c7",	x"068c0603",	x"1003102e",	x"060c0624",	
					x"062a066c",	x"065a0645",	x"065f066f",	x"0662065b",	
					x"06680663",	x"0666066a",	x"066b0652",	x"066a0684",	
					x"06a20690",	x"0692068e",	x"0698068f",	x"0694067d",	
					x"0694068b",	x"06880696",	x"06aa0662",	x"067b0661",	
					x"068b0683",	x"067f06ad",	x"06b0065f",	x"06560676",	
					x"067b0693",	x"06950675",	x"0685065a",	x"067c068f",	
					x"069106a4",	x"06a106b7",	x"069906a3",	x"069d06a2",	
					x"069a06a5",	x"068f069b",	x"06850631",	x"1003202e",	
					x"063e0626",	x"0631066c",	x"062a064b",	x"0652064a",	
					x"06640656",	x"06710651",	x"064f0655",	x"0670063c",	
					x"066f0660",	x"06780645",	x"065c0666",	x"06700673",	
					x"06780680",	x"068e066b",	x"0691067b",	x"06680628",	
					x"06530661",	x"065a066d",	x"065c0673",	x"0682067e",	
					x"068d0698",	x"06840699",	x"06800691",	x"067e0662",	
					x"0685066d",	x"06840672",	x"06780684",	x"067a069b",	
					x"0684067d",	x"06820688",	x"0677068a",	x"06670635",	
					x"1003302e",	x"05ff0644",	x"062f0637",	x"06110645",	
					x"0621064e",	x"064b0668",	x"06500653",	x"06340680",	
					x"06640653",	x"063b0650",	x"066a0670",	x"065f0664",	
					x"065c0679",	x"066d0683",	x"0679066d",	x"06690669",	
					x"064a0641",	x"06480668",	x"066d067b",	x"06730677",	
					x"067f067d",	x"067a0683",	x"0668067e",	x"0687067b",	
					x"066a066b",	x"06650686",	x"06630688",	x"066e06a3",	
					x"069306a8",	x"068c06a8",	x"0694069a",	x"066b0693",	
					x"06730626",	x"000a0004",	x"feb5dae6",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1004402e",	x"060c064a",	x"06240661",	
					x"0647065f",	x"064f067e",	x"06670681",	x"0680067e",	
					x"06860688",	x"067c067d",	x"066d0696",	x"067e068c",	
					x"06770696",	x"06980689",	x"069006a8",	x"06aa06a7",	
					x"06a7069a",	x"06a30668",	x"067306aa",	x"06ad06a5",	
					x"069406b3",	x"06cb06cd",	x"06ca069c",	x"06a306cd",	
					x"06b306c6",	x"06b0069f",	x"06a706c0",	x"06c306e8",	
					x"06d906d2",	x"06d206dd",	x"06bd06ce",	x"06d006d5",	
					x"06b606cb",	x"06bb0697",	x"1004502e",	x"0661067f",	
					x"06730699",	x"06650696",	x"069906b6",	x"067f06bc",	
					x"069c06d7",	x"06ba06bd",	x"06b606c0",	x"069c06dc",	
					x"06d106d8",	x"06bd06c2",	x"06cf06d3",	x"06b806d9",	
					x"06d006c7",	x"06b606c3",	x"06ae0697",	x"068b06d5",	
					x"06b206e1",	x"06d806dd",	x"06ca06e7",	x"06ca06eb",	
					x"06cf06ed",	x"06df06fd",	x"06cd06c9",	x"06ca06df",	
					x"06b7070f",	x"06d906ff",	x"06e60700",	x"06d606fe",	
					x"06e10703",	x"06df06f7",	x"06ec0688",	x"1004602e",	
					x"0654069d",	x"068306ae",	x"069b06b7",	x"068806c9",	
					x"06b006d5",	x"069f06ce",	x"06a206c9",	x"06b106b9",	
					x"069b06d5",	x"06c306f6",	x"06c70715",	x"06fc0712",	
					x"06ea070f",	x"06db0701",	x"06c50710",	x"06ef06de",	
					x"06ee070f",	x"070b0701",	x"06d80710",	x"06e80714",	
					x"06e90722",	x"07240710",	x"06ec0714",	x"07010713",	
					x"06f50728",	x"0704072b",	x"07030731",	x"07050730",	
					x"06e70747",	x"0729073e",	x"0708071e",	x"06fa06ba",	
					x"1004702e",	x"069e06d5",	x"069d0702",	x"06c406e6",	
					x"06c4071e",	x"06db06ee",	x"06d906e1",	x"06de073a",	
					x"06d6070d",	x"070e0741",	x"071c0743",	x"071b0747",	
					x"0731077e",	x"0737074c",	x"074c074e",	x"07380739",	
					x"0741073f",	x"071c0729",	x"074d0767",	x"0731076c",	
					x"07440780",	x"07600799",	x"07610776",	x"07570791",	
					x"076b0748",	x"072d0767",	x"0767077a",	x"078507aa",	
					x"077c07c7",	x"0782079a",	x"078607a4",	x"077f0782",	
					x"07760712",	x"000a0004",	x"2e431739",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2005002e",	x"070c071e",	x"071b0712",	
					x"06f706ee",	x"07100740",	x"07340754",	x"073d0745",	
					x"074d0729",	x"072d0719",	x"0747071d",	x"07380751",	
					x"07500764",	x"07950797",	x"0787075f",	x"07650787",	
					x"07900745",	x"0757072b",	x"073f073c",	x"075c0750",	
					x"074c0746",	x"07670784",	x"07650742",	x"07620765",	
					x"07780769",	x"07720738",	x"07520759",	x"07460761",	
					x"076d0763",	x"0780076f",	x"0762074d",	x"074c0765",	
					x"0756076a",	x"073606e4",	x"2005102e",	x"06e406e5",	
					x"06cd06ff",	x"06f7072c",	x"072d072f",	x"07550701",	
					x"072c074c",	x"0738072c",	x"0743071e",	x"07440751",	
					x"07410741",	x"07590759",	x"076d0795",	x"07720740",	
					x"075d074e",	x"0754074f",	x"0742070e",	x"074b0739",	
					x"0747074c",	x"074b0737",	x"0739073c",	x"0727074b",	
					x"07720795",	x"07720763",	x"07680730",	x"075a0753",	
					x"07560743",	x"074f076f",	x"0768076d",	x"07650762",	
					x"0762076a",	x"076d0755",	x"076406f6",	x"2005202e",	
					x"070306ed",	x"06ed06d4",	x"06ea06d6",	x"06f806f3",	
					x"0709072e",	x"074d0721",	x"07260726",	x"0750071b",	
					x"073d0711",	x"073f0721",	x"074f074d",	x"07520757",	
					x"075e0762",	x"07690749",	x"0747075b",	x"074e06d8",	
					x"07240741",	x"0757074a",	x"071c073b",	x"07380731",	
					x"0721072e",	x"07260737",	x"07390746",	x"0743070d",	
					x"07380740",	x"07540767",	x"07590759",	x"075b075e",	
					x"07410755",	x"073d0750",	x"07440754",	x"074b06f9",	
					x"2005302e",	x"06da06f4",	x"06e106fe",	x"06fd06ff",	
					x"06fe071c",	x"0719071d",	x"07060730",	x"0710071f",	
					x"073206f4",	x"07030718",	x"07280718",	x"071a0737",	
					x"0729074c",	x"07260730",	x"07260730",	x"071b072d",	
					x"06f606f2",	x"06fd071c",	x"07330734",	x"0743074e",	
					x"075e0757",	x"07410747",	x"07470751",	x"073d073d",	
					x"073d074a",	x"073c073e",	x"073a0756",	x"073e0768",	
					x"072f076a",	x"073c0752",	x"073c0759",	x"073a0763",	
					x"073e070f",	x"000a0004",	x"a2983cee",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2006402e",	x"06e70713",	x"07170711",	
					x"071d0747",	x"071a0747",	x"07390733",	x"07480743",	
					x"074b074d",	x"07640737",	x"07460745",	x"075b0763",	
					x"0769074b",	x"0765076c",	x"074e076f",	x"0763076d",	
					x"07860779",	x"074c072a",	x"075b0760",	x"075c075f",	
					x"07680778",	x"0799077f",	x"07700777",	x"0780077d",	
					x"07830792",	x"079f0772",	x"0783079b",	x"078e0787",	
					x"07840798",	x"079c07c5",	x"07a207b7",	x"07a707bd",	
					x"07a007b4",	x"0797072b",	x"2006502e",	x"073e0753",	
					x"0731074f",	x"071e0763",	x"07610783",	x"07850783",	
					x"07770787",	x"076d0791",	x"0764079a",	x"0799079b",	
					x"078807ae",	x"078b07a2",	x"07a707a1",	x"079707b3",	
					x"079e07ab",	x"07ae07a7",	x"0776077c",	x"075807ab",	
					x"078d07b7",	x"078e07ba",	x"078907ea",	x"079007da",	
					x"07a207cc",	x"079107d8",	x"07960794",	x"077d07c0",	
					x"079a07c4",	x"07a407e0",	x"07a9080a",	x"07a407e1",	
					x"07a507dd",	x"07ae07c0",	x"078a074a",	x"2006602e",	
					x"073c0771",	x"071b078a",	x"07800785",	x"07720798",	
					x"07570796",	x"0759079d",	x"07a5078a",	x"076e07ab",	
					x"077a079a",	x"077707d2",	x"07a507ce",	x"07c407f4",	
					x"07b407ea",	x"07c307e7",	x"07b807d1",	x"07cb07ab",	
					x"078807e1",	x"07d807e0",	x"07c307e9",	x"07d607f7",	
					x"07be07d0",	x"07d707ec",	x"07c407e4",	x"07d507f7",	
					x"07b4080c",	x"07d6080f",	x"07d6080b",	x"07ef0808",	
					x"080a07fb",	x"07ea080e",	x"07b6080a",	x"07d30771",	
					x"2006702e",	x"07410782",	x"075a07c6",	x"078907a9",	
					x"07a30846",	x"07a007e8",	x"07df07ed",	x"07ec07f2",	
					x"07e307e4",	x"07e30826",	x"081b082c",	x"080c082b",	
					x"082f0877",	x"0811084f",	x"07f10854",	x"07f90832",	
					x"08220810",	x"080a0852",	x"08310859",	x"081d0869",	
					x"0814085c",	x"08290858",	x"082b0862",	x"0831086b",	
					x"08580856",	x"08530861",	x"085d086d",	x"084d0893",	
					x"086508ad",	x"086a08be",	x"08630896",	x"085d0867",	
					x"086406d8",	x"000a0004",	x"d87281e2",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3007002e",	x"06c206f2",	x"06e7070c",	
					x"071406dd",	x"070906fe",	x"070106f5",	x"070f072c",	
					x"0733071e",	x"070e06dc",	x"070e0736",	x"071f073d",	
					x"073e0743",	x"07450756",	x"075c074b",	x"0732071c",	
					x"0723070e",	x"07330702",	x"072a072a",	x"0732073f",	
					x"071e0729",	x"0718075d",	x"073f072f",	x"073b0761",	
					x"076a072f",	x"07300702",	x"07330713",	x"07230714",	
					x"07290741",	x"074e0743",	x"073f073f",	x"074a0757",	
					x"07420730",	x"071706f3",	x"3007102e",	x"06d606d3",	
					x"06fc06e8",	x"06d906d9",	x"06d306ec",	x"06e906e7",	
					x"07040703",	x"071206f6",	x"070306f9",	x"070c071a",	
					x"072a0715",	x"072e0709",	x"07580706",	x"07180707",	
					x"06f90732",	x"0720072f",	x"073b070b",	x"072a0702",	
					x"07060700",	x"0700070a",	x"07380735",	x"072c0722",	
					x"0728073f",	x"07330747",	x"072606f1",	x"07200716",	
					x"070f0726",	x"07420727",	x"07370745",	x"073d0736",	
					x"072b0740",	x"073f0741",	x"073806d5",	x"3007202e",	
					x"06fb06ec",	x"070006f1",	x"070b06f1",	x"070a06e4",	
					x"071d06dd",	x"06f7071c",	x"073e0716",	x"071606cb",	
					x"06fb0702",	x"07210706",	x"07190708",	x"07080709",	
					x"07190715",	x"071d071e",	x"07060714",	x"06f706d9",	
					x"07050704",	x"06f40709",	x"070f070e",	x"070d070e",	
					x"0700071a",	x"071b0725",	x"0722072a",	x"070c06f6",	
					x"070006dd",	x"06f20721",	x"07050702",	x"0716071a",	
					x"072b0711",	x"0713072b",	x"07150736",	x"071f06cd",	
					x"3007302e",	x"06aa06cf",	x"06c506dc",	x"06d006d8",	
					x"06f506ef",	x"06c306e3",	x"06d506d3",	x"06d306d4",	
					x"06d806cb",	x"06e206fb",	x"06f106f3",	x"06e70703",	
					x"07100703",	x"06f90723",	x"070a070c",	x"07100710",	
					x"070d06e4",	x"06de06fb",	x"06f006f6",	x"06e50707",	
					x"0718070c",	x"070e0724",	x"072d0725",	x"07150716",	
					x"07090708",	x"070d0712",	x"072706fa",	x"06e10709",	
					x"07100746",	x"070d0739",	x"07280746",	x"06fd071d",	
					x"070706e7",	x"000a0004",	x"ccf72704",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3008402e",	x"06bb06e1",	x"06d406cc",	
					x"06ea06ef",	x"070506d4",	x"06ee06ee",	x"06e50707",	
					x"070f0711",	x"070b06eb",	x"07200721",	x"072b0702",	
					x"0712072e",	x"0736073a",	x"07350732",	x"072c0740",	
					x"0747071c",	x"07070706",	x"0716072d",	x"07220721",	
					x"071e073d",	x"07320747",	x"072c075c",	x"07480757",	
					x"073d0761",	x"07430708",	x"07420745",	x"073f0751",	
					x"0758075b",	x"076c0763",	x"074f0769",	x"0769077f",	
					x"07560766",	x"075b0710",	x"3008502e",	x"06ec0703",	
					x"06f2072f",	x"06fb0730",	x"07280738",	x"070a0738",	
					x"071c070f",	x"072f074e",	x"07560753",	x"07290757",	
					x"0768075e",	x"077c0753",	x"075d076b",	x"07550777",	
					x"07660773",	x"07640763",	x"0748074b",	x"071a0751",	
					x"072a075b",	x"074b076a",	x"076807ae",	x"078a0792",	
					x"0768079b",	x"07780799",	x"077a0766",	x"07480796",	
					x"076f0777",	x"075f0793",	x"0772079d",	x"076b07a3",	
					x"078307a4",	x"0768078b",	x"0760072b",	x"3008602e",	
					x"07180736",	x"071d072f",	x"074c072c",	x"070d071c",	
					x"07300751",	x"07660746",	x"07510768",	x"07540762",	
					x"07650791",	x"07750791",	x"0783078d",	x"07860797",	
					x"07720791",	x"077f0794",	x"07830792",	x"07800754",	
					x"07650783",	x"079c0796",	x"078d07ad",	x"078307d6",	
					x"07af07c6",	x"07b207c3",	x"078807b4",	x"079a07a6",	
					x"07a307c5",	x"07ac0796",	x"076c07c7",	x"07aa07f7",	
					x"07c807e9",	x"07ce07e8",	x"07bf07cf",	x"07a80755",	
					x"3008702e",	x"0735078c",	x"07740785",	x"07560759",	
					x"074807aa",	x"078e0780",	x"0779078e",	x"077e07a7",	
					x"07a507ac",	x"07b107e1",	x"07c507e9",	x"07bb07f4",	
					x"07bb07f6",	x"07c30813",	x"080c07fc",	x"07f607f7",	
					x"07fd07dd",	x"07dd07fd",	x"07fd0806",	x"07ea080a",	
					x"07e30832",	x"07fb0812",	x"083e083c",	x"081b0805",	
					x"08180817",	x"0831080b",	x"07ce082a",	x"07f1082e",	
					x"082c0880",	x"082f0878",	x"084a0877",	x"08400832",	
					x"081606cc",	x"000a0004",	x"fd3060dc",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0009002f",	x"06d906d3",	x"06f406fa",	
					x"06fd06c7",	x"06d106e3",	x"06cf06e6",	x"06d3069a",	
					x"06b30691",	x"0684066e",	x"0694069f",	x"06b906c5",	
					x"06c406bf",	x"06cf06c5",	x"06cf06de",	x"07080715",	
					x"06f90713",	x"06e706ad",	x"06c906d0",	x"06c506ca",	
					x"06d106df",	x"06f606e8",	x"06c606f2",	x"06f90708",	
					x"070f0710",	x"06e906a7",	x"06cb06d8",	x"06c106ea",	
					x"06c506f7",	x"06f406e7",	x"06d90701",	x"06f90742",	
					x"0708072d",	x"06f506bb",	x"0009102f",	x"06e306c4",	
					x"06b106ed",	x"06ba06a8",	x"069e06ce",	x"06a4069f",	
					x"06c606a1",	x"0699066f",	x"06a40667",	x"065506a3",	
					x"06a906c5",	x"069006be",	x"06cb06cf",	x"06d706e2",	
					x"06e406fb",	x"06ec06f5",	x"06e106ad",	x"06bf06a5",	
					x"06fc06d4",	x"06c206d2",	x"06ec06e1",	x"06ef06d4",	
					x"06e806c1",	x"06be06cb",	x"06b806b9",	x"06d706d4",	
					x"06e906c6",	x"06db06d9",	x"06df06e4",	x"06dd0708",	
					x"07000720",	x"06f70713",	x"070d069e",	x"0009202f",	
					x"069f06ad",	x"069c068a",	x"068006b8",	x"06a40696",	
					x"06710695",	x"06a50674",	x"06990677",	x"06830622",	
					x"0662068c",	x"06ab06bd",	x"06a906c2",	x"06cb06c9",	
					x"06ca06dd",	x"06ea06e5",	x"06d506db",	x"06d106c6",	
					x"06b406b0",	x"06b806d1",	x"06d206cb",	x"06e706d8",	
					x"06cb06dd",	x"06d906d8",	x"06c706f0",	x"06ee06b7",	
					x"06f306d7",	x"06b806d4",	x"06c206cc",	x"06ce06c9",	
					x"06c106f8",	x"06e606fe",	x"06e40702",	x"06dd069c",	
					x"0009302f",	x"065e06b6",	x"06a30698",	x"068a06a0",	
					x"0673069a",	x"067e06c7",	x"06a106a9",	x"06a00697",	
					x"06960682",	x"065606a9",	x"068a06b2",	x"06a906ce",	
					x"069506e8",	x"06c606e8",	x"06c606cd",	x"06d106d7",	
					x"06c70697",	x"06a406c4",	x"06af06ce",	x"06bb06d0",	
					x"06d006e3",	x"06ce06e9",	x"06ec06e2",	x"06d20714",	
					x"06cf06a9",	x"06cc06f5",	x"06d506ea",	x"06ae06f3",	
					x"06d80711",	x"06d30734",	x"06e5071e",	x"06fc0728",	
					x"06e806b0",	x"000a0004",	x"e6e105fd",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"000a402f",	x"069e06c4",	x"06a206cc",	
					x"068a06e1",	x"06b106f0",	x"06ad06c2",	x"069f06ce",	
					x"069306b8",	x"06a50688",	x"067606f6",	x"06be06ef",	
					x"06bd0728",	x"06d80731",	x"06e10709",	x"06f8070d",	
					x"07090714",	x"06f706ed",	x"06f70723",	x"0706071d",	
					x"06f7071f",	x"07030734",	x"07100732",	x"07220730",	
					x"07210742",	x"0700070f",	x"07050744",	x"071a073b",	
					x"06dc0737",	x"072c075d",	x"071a0763",	x"071f075e",	
					x"07130747",	x"071106e2",	x"000a502f",	x"06dd0703",	
					x"06df0717",	x"06e206f8",	x"06dd0707",	x"06e306fd",	
					x"06e70710",	x"06b7070f",	x"06ce06de",	x"06ce0737",	
					x"06d80724",	x"06c0073c",	x"070d0745",	x"071a0748",	
					x"0742074c",	x"07040740",	x"07180734",	x"06ef0750",	
					x"071e0763",	x"06eb074e",	x"07210759",	x"071f0773",	
					x"073d076b",	x"073f0756",	x"07100745",	x"07120781",	
					x"072c0776",	x"071f0778",	x"071f0787",	x"072f0791",	
					x"0752079e",	x"074b0783",	x"073c06d5",	x"000a602f",	
					x"06b70709",	x"06df06fd",	x"06e4073f",	x"06fa071c",	
					x"06f30705",	x"06d70704",	x"06c70703",	x"06f306fc",	
					x"06c30723",	x"06f4074a",	x"0728075d",	x"07200773",	
					x"0737077c",	x"07400782",	x"074e077d",	x"07400756",	
					x"072e079a",	x"07440791",	x"0745079d",	x"075807a0",	
					x"074e0780",	x"07670794",	x"074a07a0",	x"077c0765",	
					x"07540790",	x"075107c0",	x"077707b1",	x"07600813",	
					x"076907ea",	x"07a607c6",	x"078507cf",	x"07890739",	
					x"000a702f",	x"06f8073a",	x"07070757",	x"06f90735",	
					x"07070767",	x"0713074a",	x"06fb077a",	x"0721074a",	
					x"07100721",	x"06e90785",	x"073907a7",	x"075907dc",	
					x"074f07e4",	x"077107d4",	x"078507cc",	x"079607ec",	
					x"078f0782",	x"078107e0",	x"07a207dd",	x"079a07ed",	
					x"078f07f1",	x"077907fb",	x"07d307e9",	x"0793080c",	
					x"07bd07b1",	x"079307ed",	x"07bf0805",	x"07c0081e",	
					x"07be0829",	x"07d5082a",	x"07eb083a",	x"07ff081a",	
					x"07d50683",	x"000a0004",	x"16124e38",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"100b002f",	x"067e069d",	x"069306bd",	
					x"06ab0694",	x"06770663",	x"0645066b",	x"064c0670",	
					x"063b065f",	x"0637064e",	x"06690675",	x"069c0673",	
					x"067b0691",	x"06ab0685",	x"068e06a9",	x"06c606a6",	
					x"069e069c",	x"06ba066f",	x"0681068d",	x"06a406b9",	
					x"067d0685",	x"068f0699",	x"068f06a4",	x"069906a1",	
					x"06a70687",	x"06a2066c",	x"068406a4",	x"06a1069c",	
					x"06890684",	x"066706a9",	x"06b706b3",	x"069a06ba",	
					x"069406b3",	x"06990670",	x"100b102f",	x"0655067a",	
					x"06610688",	x"0686064d",	x"06580652",	x"061e0636",	
					x"06210633",	x"062b0624",	x"06750631",	x"0628064e",	
					x"0640067c",	x"066106bc",	x"06880694",	x"06870698",	
					x"069f0687",	x"068b068d",	x"069a0649",	x"06580674",	
					x"06660668",	x"0683068f",	x"06a3067e",	x"066e06a2",	
					x"06a90693",	x"06a006a5",	x"06940657",	x"066b0687",	
					x"069b06a2",	x"069706b4",	x"06ac06b7",	x"06af06c8",	
					x"06b706c3",	x"06b706a9",	x"06a20657",	x"100b202f",	
					x"065f0665",	x"066b0680",	x"06550653",	x"06400652",	
					x"06470625",	x"06380645",	x"063f0629",	x"0642061a",	
					x"063e0632",	x"064e0659",	x"066b0662",	x"0686067d",	
					x"069c0688",	x"068a0698",	x"067c0681",	x"067b0658",	
					x"0652066c",	x"0676068b",	x"068b067a",	x"06750679",	
					x"06760682",	x"0681068b",	x"06670686",	x"06870669",	
					x"068c0669",	x"06800684",	x"06730685",	x"067e068c",	
					x"066c0690",	x"068c069c",	x"0687069b",	x"0675066a",	
					x"100b302f",	x"065a0663",	x"06360662",	x"06320663",	
					x"06310641",	x"062a063f",	x"0620063e",	x"06290644",	
					x"064a0639",	x"06280622",	x"06400663",	x"063d0676",	
					x"0660069d",	x"0672068b",	x"067306a2",	x"0687068f",	
					x"065a0669",	x"065c0678",	x"066e067d",	x"06620678",	
					x"06800684",	x"06810696",	x"068106a4",	x"0685068b",	
					x"06780693",	x"067d0694",	x"067206a2",	x"06680693",	
					x"067c0694",	x"067906b0",	x"068306c0",	x"068206ab",	
					x"068b0667",	x"000a0004",	x"fe3bde00",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"100c402f",	x"0630067b",	x"065e0690",	
					x"0659066f",	x"06700672",	x"06540663",	x"0656066e",	
					x"063e0659",	x"065c066e",	x"06350679",	x"063f068b",	
					x"067806b1",	x"069106be",	x"06a106c0",	x"06a606cf",	
					x"06a506a7",	x"068006ae",	x"069706d3",	x"06be06d2",	
					x"06b606d0",	x"06d006d5",	x"06cc06ca",	x"06bb06df",	
					x"06ce06be",	x"06b406b9",	x"06c006d5",	x"06ac06d3",	
					x"06b806df",	x"06c406eb",	x"06c60700",	x"06e406f0",	
					x"06bf0701",	x"06dc0698",	x"100c502f",	x"06850688",	
					x"06780688",	x"067a0697",	x"068506a5",	x"068506a6",	
					x"068306c0",	x"06b106b0",	x"06820694",	x"068d06e1",	
					x"06aa06cb",	x"068406d1",	x"06cc06fb",	x"06b40707",	
					x"06c506ea",	x"06bb06f7",	x"06cd06c7",	x"069c06d3",	
					x"06b90702",	x"06bc0713",	x"06da0713",	x"06d3070c",	
					x"06e60701",	x"06e60705",	x"06d606f6",	x"06d106f2",	
					x"06c0070f",	x"06db072d",	x"06dc0731",	x"06ed072f",	
					x"06fe072e",	x"06f50715",	x"06ea06ae",	x"100c602f",	
					x"068d06c3",	x"067706d5",	x"068206a9",	x"067006a5",	
					x"067a06cd",	x"066a06a9",	x"067106a6",	x"068006a9",	
					x"069306b7",	x"069b06c4",	x"0699070f",	x"06e90722",	
					x"06f2071f",	x"06fe0710",	x"06d906ff",	x"06d306e2",	
					x"06c5072d",	x"07260717",	x"06ff072c",	x"07080736",	
					x"06f5073b",	x"07080742",	x"071c0741",	x"06fe072e",	
					x"0700072f",	x"07090724",	x"06fb074c",	x"070f073a",	
					x"07100762",	x"072a074e",	x"072b0737",	x"071d06f8",	
					x"100c702f",	x"068606d4",	x"069b06d0",	x"06b506f1",	
					x"06c506d9",	x"066f06e3",	x"06c506f2",	x"06b006e3",	
					x"06ce06c3",	x"069e072d",	x"07020726",	x"07180744",	
					x"0728075f",	x"071a0762",	x"0759077e",	x"07120735",	
					x"071b0728",	x"06ee0773",	x"07260766",	x"0725077b",	
					x"076d0795",	x"075007a2",	x"074f0791",	x"0747078e",	
					x"075a075a",	x"074f0798",	x"076a07ad",	x"07530798",	
					x"077307ca",	x"078707c3",	x"079b07b7",	x"079f07ae",	
					x"07710703",	x"000a0004",	x"2bff1d1a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"200d002f",	x"0716072c",	x"07600729",	
					x"0720070a",	x"07210730",	x"07250728",	x"06f50713",	
					x"07090738",	x"074d071e",	x"07520771",	x"07680773",	
					x"0778075d",	x"07770762",	x"07640766",	x"07730799",	
					x"077d0757",	x"072d0716",	x"07390751",	x"07860746",	
					x"07610745",	x"07670756",	x"07600759",	x"0764075c",	
					x"07680771",	x"076d0748",	x"076c076c",	x"077807a4",	
					x"07810787",	x"076a0759",	x"0766076c",	x"07610779",	
					x"07640779",	x"075f06ec",	x"200d102f",	x"070a0719",	
					x"07100738",	x"07410702",	x"071b06fd",	x"06db06f4",	
					x"07150713",	x"0735071b",	x"072906e4",	x"0711073a",	
					x"0731074f",	x"07720760",	x"076c075e",	x"074b0754",	
					x"07600764",	x"076a075d",	x"0759070b",	x"070a071f",	
					x"072f073f",	x"0745075b",	x"075c0768",	x"075a0730",	
					x"0750076e",	x"074a0758",	x"07670749",	x"0760075a",	
					x"075b075f",	x"075e078a",	x"07760763",	x"075d0766",	
					x"07550770",	x"07520764",	x"075a06fe",	x"200d202f",	
					x"07200714",	x"071306fa",	x"07060705",	x"071e06fa",	
					x"06f006f9",	x"071f06fa",	x"07160744",	x"073406e8",	
					x"070c0721",	x"073c0757",	x"07460748",	x"074d0754",	
					x"073d073d",	x"07460750",	x"0746074e",	x"07360712",	
					x"0706073e",	x"0762074a",	x"073a0734",	x"07390731",	
					x"073e073a",	x"07370754",	x"0750074d",	x"074e0748",	
					x"0757075c",	x"07460756",	x"073d075a",	x"0754074c",	
					x"07260754",	x"0749074a",	x"073c075f",	x"075506cc",	
					x"200d302f",	x"06b7070c",	x"06ff071d",	x"06fb070b",	
					x"06fb06ef",	x"06d006f1",	x"06d3071d",	x"06e3070f",	
					x"07070708",	x"06f7072f",	x"07300760",	x"07440754",	
					x"07460748",	x"07410749",	x"07500744",	x"072f0743",	
					x"07180713",	x"07220755",	x"074c073e",	x"07400744",	
					x"07460763",	x"074c077f",	x"075b0795",	x"0750076d",	
					x"075a076a",	x"074a0777",	x"0748076b",	x"074f077e",	
					x"073c0777",	x"0748077d",	x"07690784",	x"07470783",	
					x"074f070d",	x"000a0004",	x"a37240dd",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"200e402f",	x"07070749",	x"070d0729",	
					x"06f20710",	x"06e40715",	x"06f7072a",	x"072c072d",	
					x"07250773",	x"0739074f",	x"075b0769",	x"07790776",	
					x"07600761",	x"076d076c",	x"07650786",	x"076c0775",	
					x"07750771",	x"075f0773",	x"0759078b",	x"07830780",	
					x"0771079a",	x"077507b4",	x"075d07b6",	x"079307ae",	
					x"078d07bb",	x"07ae0792",	x"078f07c1",	x"07b207b4",	
					x"07a007c7",	x"07a107af",	x"079007c2",	x"07b207d8",	
					x"07a807d7",	x"07970769",	x"200e502f",	x"0739077f",	
					x"07710794",	x"0740077d",	x"07560775",	x"07190758",	
					x"072c079a",	x"0777078b",	x"073c0788",	x"079507a1",	
					x"076b07c2",	x"079107d6",	x"07a207c9",	x"079c07b4",	
					x"079a07a2",	x"07a307d7",	x"078a0798",	x"077b07cf",	
					x"07c107d1",	x"079607dc",	x"07ab07ea",	x"07a407e2",	
					x"07a707f3",	x"07a707fe",	x"07aa07c7",	x"0799080b",	
					x"07a907d2",	x"07a607e9",	x"07a807f9",	x"07a60814",	
					x"07c6080e",	x"07ba0801",	x"07a4075d",	x"200e602f",	
					x"07380786",	x"076b0782",	x"0768077e",	x"074e079b",	
					x"0764078c",	x"0765077d",	x"0760078b",	x"07690797",	
					x"075d07fe",	x"079c0802",	x"07aa0813",	x"07cf0819",	
					x"07aa07ec",	x"07b407d6",	x"07bd07ce",	x"07c307d2",	
					x"07b207e4",	x"07c0080c",	x"07b50821",	x"07d3080c",	
					x"07c40833",	x"0812083b",	x"07e6082b",	x"07bd07fc",	
					x"07d8082a",	x"07d0081e",	x"07ce085c",	x"07e7082b",	
					x"07e3084f",	x"08110834",	x"07e70841",	x"07d807b3",	
					x"200e702f",	x"076a07d8",	x"07700789",	x"076e07c4",	
					x"077d07e9",	x"078607bd",	x"076807d4",	x"077507ec",	
					x"07aa07fd",	x"07f10845",	x"0804084b",	x"08030862",	
					x"08110853",	x"08070850",	x"08010876",	x"0839083f",	
					x"08010847",	x"08120849",	x"080e082c",	x"08090891",	
					x"082f0897",	x"0823088e",	x"084b0885",	x"0860088c",	
					x"0851084d",	x"0841088e",	x"085f0888",	x"085808ba",	
					x"08870899",	x"085408b0",	x"085608b0",	x"086a08ad",	
					x"08520743",	x"000a0004",	x"d8418ddf",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"300f002f",	x"071006ec",	x"070506fb",	
					x"06ee06ea",	x"06f406e2",	x"06f006e6",	x"06f306fd",	
					x"06ed0711",	x"074606fa",	x"06fd0739",	x"073a0735",	
					x"07520746",	x"0759076d",	x"075c0764",	x"0761074e",	
					x"07630728",	x"074c06f4",	x"0727072b",	x"07400733",	
					x"073c0721",	x"073a0734",	x"071b077f",	x"0763076c",	
					x"0758074f",	x"073e0707",	x"0748074c",	x"07560749",	
					x"071c0741",	x"0733074a",	x"072e073f",	x"07490779",	
					x"074f076a",	x"075306d4",	x"300f102f",	x"06d406e7",	
					x"06fe06f6",	x"06e906c3",	x"06c406c2",	x"06dd06c3",	
					x"06eb06ec",	x"06e20703",	x"06d706f0",	x"06f306ff",	
					x"07220741",	x"074b0740",	x"0760075a",	x"073b0736",	
					x"0749072a",	x"07230702",	x"070f06e5",	x"06fa06ec",	
					x"0708070b",	x"06f80732",	x"07520738",	x"0729071f",	
					x"0744071c",	x"0727074a",	x"07350716",	x"0751072e",	
					x"07540754",	x"0723073e",	x"071e0726",	x"071d072c",	
					x"073b0744",	x"073f074a",	x"076106f2",	x"300f202f",	
					x"06d606e4",	x"06d806d6",	x"06d606f2",	x"06fe06d1",	
					x"06ec06d7",	x"06e006f9",	x"06f506ac",	x"06db06a0",	
					x"06f906f2",	x"07310718",	x"07240720",	x"070a0714",	
					x"071b0713",	x"0729070e",	x"0701070a",	x"070706cb",	
					x"06ee0711",	x"0726070a",	x"06f30702",	x"070b070d",	
					x"07090725",	x"07180739",	x"073b0737",	x"07210712",	
					x"07250724",	x"0722072d",	x"071f0736",	x"07240732",	
					x"071d071b",	x"070e0726",	x"0714073e",	x"071006e1",	
					x"300f302f",	x"06c906f6",	x"06d206da",	x"06cd06c6",	
					x"06ac06cf",	x"06a706d3",	x"06c606c6",	x"06c706e2",	
					x"06c306c0",	x"06d30701",	x"070c071a",	x"06f30717",	
					x"07190726",	x"0702072d",	x"071b072e",	x"070a0706",	
					x"06f906e3",	x"06d80720",	x"071c071b",	x"06f3072b",	
					x"072b0725",	x"071b071e",	x"0719073f",	x"071e073c",	
					x"07120740",	x"07220741",	x"072e072a",	x"0700071d",	
					x"070b072b",	x"07050730",	x"07020749",	x"0701073d",	
					x"070e06f7",	x"000a0004",	x"ce0d2a9c",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3010402f",	x"06d306e6",	x"06d006e3",	
					x"06de06ee",	x"06fa06fe",	x"06f00708",	x"06ec06f9",	
					x"06f4072a",	x"071f0707",	x"06ed073d",	x"07300732",	
					x"072c0732",	x"072c074d",	x"072f0751",	x"0731074a",	
					x"07260733",	x"07010713",	x"07110754",	x"074b076d",	
					x"07440769",	x"07540776",	x"074f0776",	x"075b0775",	
					x"075d0788",	x"0759074f",	x"0760076c",	x"07630770",	
					x"075b075d",	x"0761078e",	x"07550788",	x"07650795",	
					x"075e0782",	x"074b072e",	x"3010502f",	x"06b4074e",	
					x"07070731",	x"06e30738",	x"0725074c",	x"06f10762",	
					x"07600750",	x"072a0759",	x"072c0759",	x"0755079a",	
					x"0776079d",	x"0772076e",	x"0769079e",	x"075f0794",	
					x"07730773",	x"0766076c",	x"07460753",	x"07450785",	
					x"07710780",	x"077107a7",	x"077607af",	x"079407ba",	
					x"078a07b8",	x"07a807b1",	x"077207a0",	x"077807ce",	
					x"079107b3",	x"077f0795",	x"0777079f",	x"076107ec",	
					x"078b07ca",	x"079707bf",	x"078b0759",	x"3010602f",	
					x"0717076e",	x"073c076f",	x"071e0758",	x"07010738",	
					x"0715073b",	x"07400769",	x"071f075c",	x"07370769",	
					x"074507c7",	x"075d07a2",	x"079507ac",	x"079c07bc",	
					x"079107a3",	x"079907b3",	x"078407c7",	x"078d0781",	
					x"076f07c9",	x"07a707d3",	x"078807dc",	x"07b207ef",	
					x"07ac080a",	x"07bc07de",	x"07ac07ff",	x"07ae07b7",	
					x"07a907e6",	x"07c007d2",	x"07a807ce",	x"07a607f0",	
					x"07bd080f",	x"07cc0807",	x"07c10807",	x"079c074f",	
					x"3010702f",	x"0728079a",	x"07470777",	x"074407ab",	
					x"074a0770",	x"076e07b5",	x"078407e6",	x"077307b1",	
					x"078b07ac",	x"07830812",	x"07be0811",	x"07cd081c",	
					x"07da0834",	x"07e60816",	x"07f80846",	x"080a0804",	
					x"07e307d2",	x"07c40826",	x"08060830",	x"07ef0831",	
					x"081e085d",	x"07fa0834",	x"081a0880",	x"082d086a",	
					x"0820082a",	x"08370846",	x"082c084e",	x"0826085c",	
					x"08350884",	x"08140881",	x"083e0888",	x"083b0882",	
					x"081f069f",	x"000a0004",	x"00587114",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"00110030",	x"06eb069a",	x"06820695",	
					x"067a0698",	x"067d068f",	x"067306c0",	x"06c506eb",	
					x"06f806cb",	x"06c40684",	x"06ae06e0",	x"06e006d6",	
					x"06c406c0",	x"06dc06dc",	x"06d206dc",	x"06f006df",	
					x"06dc06de",	x"06d6068d",	x"069a06cd",	x"070a06eb",	
					x"06d506b8",	x"06de06c4",	x"06a406dc",	x"06e106ef",	
					x"06ec06c3",	x"06c806bb",	x"06c506da",	x"06e706e8",	
					x"06d806f3",	x"06f606f7",	x"06d706d2",	x"06c006da",	
					x"06c206fd",	x"06f206a6",	x"00111030",	x"06b40667",	
					x"069006a5",	x"06b70673",	x"069906a5",	x"069f06a3",	
					x"06a606c9",	x"06c50696",	x"06c406b0",	x"06a006b4",	
					x"06bc06bf",	x"06e406bc",	x"06ef06c0",	x"06d606ba",	
					x"06cd06c2",	x"06db06df",	x"06d0067e",	x"069a06b9",	
					x"06c106de",	x"06e206ca",	x"06d006c4",	x"06cf06c2",	
					x"06df06d2",	x"06e106d0",	x"06d106b6",	x"06c106cb",	
					x"06bd06db",	x"06dd06fa",	x"070706fd",	x"06ea06eb",	
					x"06da06f9",	x"070906ee",	x"06f90676",	x"00112030",	
					x"06ba0673",	x"0693069c",	x"067d066c",	x"0687068a",	
					x"06a3068e",	x"06b2069f",	x"06a50699",	x"06c10686",	
					x"06ca06d2",	x"06df06d1",	x"06db06d2",	x"06d806bc",	
					x"06b706ba",	x"06bf06cd",	x"06be06ab",	x"06ac0687",	
					x"06a606f0",	x"06c706c8",	x"06d006be",	x"06cd06ba",	
					x"06b306e4",	x"06c206d9",	x"06d406d5",	x"06cc069d",	
					x"06ab06d9",	x"06ce06da",	x"06c806cd",	x"06d506d3",	
					x"06cf06eb",	x"06ee06e8",	x"06d406e0",	x"06be066d",	
					x"00113030",	x"06750676",	x"065f0690",	x"069206ad",	
					x"0682068b",	x"068806a6",	x"06a506ba",	x"069b06b2",	
					x"0695068f",	x"069906d7",	x"06c506b3",	x"06a006b6",	
					x"06a806b9",	x"06a106c9",	x"06b106b2",	x"069506c6",	
					x"06b60689",	x"06a406c6",	x"06b606cf",	x"06a006cf",	
					x"06d706f5",	x"06d106f7",	x"06cb06d5",	x"06b306cf",	
					x"06cc0696",	x"06aa06e4",	x"06d5070f",	x"06d706f2",	
					x"06dc06de",	x"06be0700",	x"06ca06ec",	x"06d10707",	
					x"06e00699",	x"000a0004",	x"e4a10026",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"00124030",	x"068f06af",	x"06ad06a4",	
					x"0692069a",	x"069f06d1",	x"06b306cf",	x"06ae06d0",	
					x"06ec06b9",	x"06a906b8",	x"06c106f0",	x"06e106f9",	
					x"06ce06fd",	x"06f20710",	x"06e006e8",	x"06ec06e9",	
					x"06f006ff",	x"06f006d4",	x"06e1070c",	x"0710071d",	
					x"0708070e",	x"07000717",	x"06fa071a",	x"071c0715",	
					x"070f070a",	x"06f70709",	x"07130727",	x"071f0729",	
					x"07160740",	x"07350744",	x"07130743",	x"071b0751",	
					x"07090746",	x"071906d0",	x"00125030",	x"06ee06dc",	
					x"06bf0700",	x"06f506e0",	x"06e006f7",	x"06ea0717",	
					x"06e5072b",	x"0709073c",	x"07250714",	x"06fa0738",	
					x"0719073c",	x"071a0749",	x"07360744",	x"071a0739",	
					x"070f0734",	x"06f50725",	x"07000726",	x"06ff0752",	
					x"0729072c",	x"0703073a",	x"07170743",	x"071b074f",	
					x"073b074f",	x"071c0760",	x"073d0751",	x"07050764",	
					x"0740076f",	x"0742076d",	x"07300781",	x"07300780",	
					x"073c0775",	x"071e0769",	x"07310704",	x"00126030",	
					x"06f60725",	x"06f70713",	x"06c30739",	x"06f30723",	
					x"06f40736",	x"07120747",	x"0708074d",	x"072a0736",	
					x"071a076d",	x"07330773",	x"07580765",	x"074d0761",	
					x"07510757",	x"07730789",	x"0757075e",	x"073b075f",	
					x"073f075b",	x"076b077a",	x"0756077c",	x"0772077f",	
					x"0748076f",	x"074a0787",	x"07440780",	x"0758077f",	
					x"0756078e",	x"077507ac",	x"077c07a1",	x"078407bf",	
					x"077007bc",	x"077807af",	x"076f07b3",	x"077c0760",	
					x"00127030",	x"075d076e",	x"0727075b",	x"07130771",	
					x"073c07ae",	x"07440779",	x"07670793",	x"0785079a",	
					x"076d0795",	x"076807c0",	x"07ab07c1",	x"07a607c4",	
					x"079507ca",	x"07a807bc",	x"079b07ce",	x"07af07c9",	
					x"07ac07c6",	x"07b907f9",	x"07c107ee",	x"07c20812",	
					x"07d907fc",	x"07db07e0",	x"07cb07f9",	x"07cc07e3",	
					x"07ef07e9",	x"07d407ff",	x"07ed081b",	x"07e70810",	
					x"08010852",	x"08110836",	x"08190835",	x"081d0822",	
					x"07fe064f",	x"000a0004",	x"220f4d6e",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"10130030",	x"06470646",	x"065c0654",	
					x"065f065c",	x"066b067b",	x"06a10683",	x"066d0683",	
					x"065e0675",	x"06670667",	x"0677067f",	x"06c10674",	
					x"067806a2",	x"06960691",	x"0696069c",	x"06ba069d",	
					x"06a30695",	x"06ad0652",	x"066e066f",	x"065e0689",	
					x"06760678",	x"0685067e",	x"06950695",	x"067e06ba",	
					x"06b2068e",	x"06a60642",	x"0655067d",	x"069506a7",	
					x"069b06a3",	x"06b8068e",	x"069b068f",	x"06a00698",	
					x"067a0694",	x"067e061e",	x"10131030",	x"0633062d",	
					x"06320641",	x"063f064c",	x"066b0671",	x"0672066d",	
					x"066f0693",	x"068a0665",	x"068c065a",	x"066e0663",	
					x"06830679",	x"067a0686",	x"06aa0691",	x"06800681",	
					x"0698068b",	x"068a067f",	x"06920667",	x"06650658",	
					x"066d0663",	x"0672068a",	x"069a0674",	x"067c0698",	
					x"06b206aa",	x"06bb068e",	x"068f0683",	x"067d0677",	
					x"06820695",	x"06aa06c3",	x"06b20698",	x"06a206ac",	
					x"0692068d",	x"06930698",	x"06a3064e",	x"10132030",	
					x"066a063b",	x"0650064e",	x"0652065b",	x"0658063a",	
					x"065b065b",	x"066b067a",	x"06630647",	x"0664063e",	
					x"06810673",	x"06870669",	x"066e0649",	x"0666067d",	
					x"067c0680",	x"0673067e",	x"067f0672",	x"06780646",	
					x"06440685",	x"066a0674",	x"064e0660",	x"06750672",	
					x"067c0699",	x"0696069e",	x"068d067a",	x"0668064d",	
					x"0667068a",	x"06890698",	x"066d068f",	x"06910693",	
					x"067a068a",	x"06770678",	x"06630685",	x"066e063e",	
					x"10133030",	x"063c0634",	x"0617063f",	x"0629065b",	
					x"06430656",	x"064f0661",	x"06570656",	x"06550675",	
					x"066d064a",	x"06380658",	x"06620652",	x"0657066c",	
					x"0665067c",	x"0656066d",	x"06700676",	x"06650666",	
					x"064e0663",	x"065e0663",	x"066e066e",	x"06770676",	
					x"067e0677",	x"0674067e",	x"066c0677",	x"0670068c",	
					x"066c0686",	x"0664069e",	x"06740693",	x"06780699",	
					x"068f069e",	x"067f0696",	x"06890695",	x"06660689",	
					x"066d064c",	x"000a0004",	x"ff74da78",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"10144030",	x"062b064f",	x"061e066c",	
					x"06400683",	x"065d0689",	x"06620681",	x"06830686",	
					x"067d0692",	x"0684067b",	x"067306a1",	x"06880694",	
					x"067d068e",	x"06920699",	x"069206a9",	x"06a106a2",	
					x"06a70698",	x"06a0067a",	x"068906ae",	x"06b406af",	
					x"06a0069b",	x"06ba06ad",	x"06bf06a2",	x"06ac06c8",	
					x"06b506ca",	x"06bc06af",	x"06ab06c2",	x"06a806cc",	
					x"06ca06c6",	x"06d806d6",	x"06be06e0",	x"06c506cc",	
					x"069b06df",	x"06bb0698",	x"10145030",	x"06960680",	
					x"066906a3",	x"067306a2",	x"06ad06b2",	x"06a606cf",	
					x"06b106d7",	x"06cb06cd",	x"06de06bc",	x"06c306ce",	
					x"06c106cf",	x"06c506db",	x"06d606de",	x"06bc06c9",	
					x"06b006c9",	x"06b306ce",	x"06be06b7",	x"06b306ce",	
					x"06c406de",	x"06cb06e8",	x"06d106fe",	x"06db06f0",	
					x"06db06f8",	x"06e506fd",	x"06df06f0",	x"06cb06f6",	
					x"06c40712",	x"06cb070b",	x"06e806f8",	x"06ce06ec",	
					x"06df0708",	x"06e406fb",	x"06e606a8",	x"10146030",	
					x"067e06bd",	x"068206cf",	x"068106b4",	x"06ad06d0",	
					x"06df06db",	x"06cb06f8",	x"06c706f5",	x"06dc06bc",	
					x"06c106fc",	x"06e4070a",	x"06c30715",	x"06fc070c",	
					x"06f20704",	x"06f106ff",	x"06db0721",	x"06da06d3",	
					x"06c90711",	x"070206f9",	x"06e6070b",	x"070b072f",	
					x"07230728",	x"071a072a",	x"070a071d",	x"07010706",	
					x"06f7073a",	x"07260731",	x"0710072d",	x"0704072d",	
					x"07160740",	x"07250746",	x"071d072a",	x"0707070b",	
					x"10147030",	x"06d90712",	x"06e30706",	x"06f5072a",	
					x"071d0729",	x"06ff0711",	x"07130722",	x"06fa071b",	
					x"071a0736",	x"072a0762",	x"074b0745",	x"072b0757",	
					x"075b0770",	x"07440775",	x"075a077c",	x"07570761",	
					x"07520762",	x"0738076e",	x"07580772",	x"07680772",	
					x"076207b5",	x"077f07b9",	x"07890799",	x"07590776",	
					x"0759075a",	x"075a07a1",	x"079b0792",	x"07a8078b",	
					x"079007c1",	x"079007bc",	x"07b707b7",	x"079a07a8",	
					x"07820709",	x"000a0004",	x"36171ce9",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"20150030",	x"07490701",	x"07030702",	
					x"070c070f",	x"07190720",	x"072c074d",	x"073f074e",	
					x"0743074f",	x"076a072d",	x"073c0729",	x"07620724",	
					x"074e0751",	x"075a0758",	x"07740769",	x"07920773",	
					x"0782074e",	x"075706f3",	x"07410734",	x"074b0755",	
					x"07530734",	x"07490752",	x"07530741",	x"07550747",	
					x"07530746",	x"075b071c",	x"071f0732",	x"0734074c",	
					x"0742074f",	x"0751076a",	x"071f073c",	x"0745077d",	
					x"0744076f",	x"075306e1",	x"20151030",	x"06ed06f6",	
					x"07060705",	x"070106fd",	x"06f20740",	x"0731072c",	
					x"073d0731",	x"073d072c",	x"074b070c",	x"07160733",	
					x"07410734",	x"07310770",	x"07850790",	x"0752075d",	
					x"0770075d",	x"07440747",	x"07460706",	x"071d0725",	
					x"074f0749",	x"075a0757",	x"075c073e",	x"0737072e",	
					x"0740077c",	x"07640769",	x"07570720",	x"0736075a",	
					x"075f076a",	x"07660763",	x"07650752",	x"074c0745",	
					x"074c0789",	x"07710763",	x"076206eb",	x"20152030",	
					x"06ec070b",	x"071206fc",	x"070d0708",	x"07420713",	
					x"072d071f",	x"07430720",	x"07320711",	x"072c06f5",	
					x"070f0705",	x"07400709",	x"07360724",	x"07300756",	
					x"0758074a",	x"074f0734",	x"07520759",	x"073406c4",	
					x"071c0727",	x"0728071b",	x"070e0727",	x"07360727",	
					x"0731072c",	x"07430767",	x"074c073c",	x"073f071f",	
					x"07310747",	x"073d0752",	x"0726073e",	x"0762074b",	
					x"0740074b",	x"07320747",	x"07310737",	x"075206d2",	
					x"20153030",	x"06cf06e7",	x"06ce06f1",	x"070006f1",	
					x"070506f6",	x"06fe0712",	x"0708072e",	x"07180708",	
					x"071906ec",	x"07040709",	x"0722072d",	x"073c0749",	
					x"07360738",	x"0727073f",	x"0751073a",	x"0715072e",	
					x"073306f2",	x"0707072c",	x"072a0730",	x"073b0739",	
					x"0738074d",	x"0740074e",	x"073d0750",	x"073a074d",	
					x"07410703",	x"07130734",	x"072c0756",	x"07320768",	
					x"07320762",	x"0738075c",	x"074f077b",	x"07380774",	
					x"0742070a",	x"000a0004",	x"a08439b8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"20164030",	x"070a0711",	x"07240714",	
					x"071e0742",	x"071e074a",	x"0730074a",	x"07610749",	
					x"07330741",	x"07440728",	x"074c0736",	x"07500761",	
					x"076e075d",	x"07600774",	x"07580783",	x"077e077e",	
					x"074d0761",	x"074b0737",	x"0756076b",	x"075d0769",	
					x"076e0778",	x"077f0794",	x"077a077e",	x"077e078d",	
					x"079b0780",	x"077f078d",	x"077c0792",	x"07910787",	
					x"077e079e",	x"079907ba",	x"079a07a5",	x"0799079e",	
					x"079207c4",	x"07a90730",	x"20165030",	x"0748074f",	
					x"07230775",	x"074e076d",	x"07640775",	x"0773079a",	
					x"07730775",	x"077e0773",	x"075b07a0",	x"07a507a8",	
					x"07a407ad",	x"0791079d",	x"079907d0",	x"07b507af",	
					x"07a807ad",	x"07aa07bc",	x"07840792",	x"076507ae",	
					x"07aa07bb",	x"079d07d9",	x"07b007c7",	x"07a707bb",	
					x"07aa07df",	x"07ac07d3",	x"07a507b5",	x"079407bb",	
					x"07a407da",	x"07a207e0",	x"07a107fb",	x"07ac07f7",	
					x"07b507ec",	x"07af07de",	x"07af0778",	x"20166030",	
					x"07510777",	x"075d076d",	x"07590771",	x"0757079c",	
					x"0779079e",	x"077c07ae",	x"078807a9",	x"079307c1",	
					x"078307e2",	x"078d07e7",	x"07c307e5",	x"07c107ff",	
					x"07b707ed",	x"07ce07f8",	x"07aa07cd",	x"07c607db",	
					x"07bf07e2",	x"07df07d8",	x"07c00804",	x"07e307fe",	
					x"07be07f8",	x"08030802",	x"07c3080c",	x"07f90800",	
					x"07ef0804",	x"07df081a",	x"07de0827",	x"0804081d",	
					x"07f80815",	x"07d7081f",	x"07e80835",	x"07f107e0",	
					x"20167030",	x"07a407bb",	x"07a807fb",	x"077e07e4",	
					x"07c70819",	x"07e80809",	x"0815081c",	x"08170810",	
					x"07ed07e7",	x"07e70838",	x"0822083f",	x"08330849",	
					x"084a0896",	x"08250863",	x"082a0855",	x"08330855",	
					x"081c0840",	x"08370843",	x"083f088d",	x"08380880",	
					x"086d0880",	x"08570874",	x"084e087f",	x"0858088a",	
					x"08560867",	x"084d0885",	x"087c088e",	x"088c08a0",	
					x"08900893",	x"087c08af",	x"089808bd",	x"088f0894",	
					x"08960710",	x"000a0004",	x"e03788bc",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"30170030",	x"06f306d2",	x"06dd06d2",	
					x"06d006d4",	x"06ec06c9",	x"070906ee",	x"06f70713",	
					x"07330717",	x"071f06f2",	x"06fa0723",	x"0729071c",	
					x"071f0717",	x"07550743",	x"070d073a",	x"0726073e",	
					x"074906f7",	x"06fe06d4",	x"06fc070f",	x"07170717",	
					x"071306f5",	x"0702072f",	x"06fe0717",	x"073b0766",	
					x"07550737",	x"071e06f3",	x"06e70710",	x"07170716",	
					x"07150722",	x"073b0727",	x"0710072c",	x"07270765",	
					x"073f0750",	x"071c06cf",	x"30171030",	x"06ea06d9",	
					x"06eb06fa",	x"06f006dc",	x"06d706e1",	x"06df06ec",	
					x"07190719",	x"071606e4",	x"06f206d8",	x"06f2070d",	
					x"07330729",	x"073c0712",	x"07430718",	x"070a071e",	
					x"0718070b",	x"0719070f",	x"073606dc",	x"06d10702",	
					x"072206e8",	x"06ee0705",	x"07420718",	x"07240707",	
					x"073d0729",	x"072e0730",	x"071c06fe",	x"06f106f6",	
					x"06fa06fb",	x"07190721",	x"0719072a",	x"07150740",	
					x"073c0739",	x"072e0734",	x"072c06ed",	x"30172030",	
					x"06ee06e6",	x"06f406eb",	x"06e606c8",	x"06da06d0",	
					x"070106d6",	x"06f906fc",	x"070406ee",	x"071a06ef",	
					x"0712070b",	x"072706f8",	x"07370712",	x"0705070b",	
					x"070a0706",	x"07180723",	x"06f806f7",	x"070406e7",	
					x"06f706ec",	x"06f306ed",	x"06d306ec",	x"06f206f6",	
					x"0706072d",	x"0734072e",	x"0727071f",	x"070a06f2",	
					x"06f806f5",	x"06f306f9",	x"06fe0708",	x"0705071c",	
					x"070e072f",	x"071d0717",	x"06f70730",	x"071206d5",	
					x"30173030",	x"06d206dc",	x"06e506e1",	x"06d206b1",	
					x"06c906db",	x"06b606e7",	x"06dc06e6",	x"06e506ec",	
					x"06d306de",	x"06e306e4",	x"071206ff",	x"06fd0722",	
					x"071c06ee",	x"06e20701",	x"06f606f7",	x"06f806f1",	
					x"06e506d0",	x"06cd06f7",	x"06f80706",	x"06ef0711",	
					x"071106f4",	x"06e20716",	x"07180728",	x"07080715",	
					x"06ee06fe",	x"06fa071d",	x"0727070f",	x"06fe0717",	
					x"07070737",	x"07100731",	x"071c0746",	x"06fa0715",	
					x"070806e5",	x"000a0004",	x"c8262260",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"30184030",	x"06ce06f1",	x"06d206f9",	
					x"06fd0709",	x"06fb06ec",	x"06e80704",	x"0708070a",	
					x"071b070a",	x"0704070f",	x"0717070e",	x"072b071a",	
					x"0711072a",	x"070f072e",	x"0718072f",	x"072a073e",	
					x"073c0729",	x"072b0715",	x"07290729",	x"0721072d",	
					x"0728072b",	x"0735073e",	x"07360751",	x"07370757",	
					x"073d075f",	x"07580710",	x"072f0743",	x"07400752",	
					x"074e075c",	x"07690788",	x"07670781",	x"07710775",	
					x"074a0769",	x"0742074b",	x"30185030",	x"0735070f",	
					x"06f90730",	x"06ef072a",	x"07260741",	x"07220757",	
					x"074f0755",	x"073b0755",	x"073b0761",	x"0756075e",	
					x"0764075c",	x"0766075a",	x"07650755",	x"07550783",	
					x"076a0766",	x"076a0764",	x"075d0760",	x"072a0756",	
					x"0748075c",	x"075f0773",	x"0770078b",	x"077407bb",	
					x"078f07a7",	x"078e078e",	x"07780779",	x"07570793",	
					x"07470783",	x"077807ae",	x"078207ac",	x"077b07be",	
					x"078307bf",	x"078f079e",	x"07760755",	x"30186030",	
					x"07230767",	x"0751074f",	x"07300742",	x"07310770",	
					x"0774076e",	x"075d075c",	x"07490761",	x"075b0773",	
					x"076a078e",	x"07790798",	x"078f079c",	x"079707a9",	
					x"078f079b",	x"079c0799",	x"077407a0",	x"0774076f",	
					x"0779078f",	x"079307ad",	x"079107ac",	x"078b07c7",	
					x"079c07c0",	x"07b307d2",	x"07b107c4",	x"07b007c4",	
					x"07a707d1",	x"07a507aa",	x"079c07cf",	x"07b407ff",	
					x"07c207da",	x"07c907e5",	x"07a407e0",	x"07bc0760",	
					x"30187030",	x"075c07a3",	x"078307a7",	x"077f07a4",	
					x"077f07b2",	x"079c07c4",	x"07bc07e4",	x"07ba07a4",	
					x"07c107b3",	x"07da0814",	x"07f807f5",	x"07f607f3",	
					x"07f3080d",	x"0805082d",	x"081e0838",	x"0807080d",	
					x"07fc07cf",	x"07cf080e",	x"07fb081e",	x"080c081c",	
					x"081f0850",	x"081f0838",	x"085a085f",	x"08540836",	
					x"08450826",	x"08470832",	x"08460863",	x"083f0866",	
					x"08500874",	x"08480892",	x"085a0885",	x"08640863",	
					x"086706b6",	x"000a0004",	x"053568b9",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"00190031",	x"06dc06c1",	x"06c206c2",	
					x"06c806d8",	x"06cf06ce",	x"06ae06b9",	x"069b0692",	
					x"0684069f",	x"06a50670",	x"067e06b4",	x"06b606ad",	
					x"06ab06b9",	x"06be06c5",	x"06c106bf",	x"06e306cc",	
					x"06d406d1",	x"06ba06a2",	x"06bb06e0",	x"06c706c3",	
					x"06c406d3",	x"06e506d0",	x"06a506f2",	x"06e50706",	
					x"07150708",	x"06ec0693",	x"069206c3",	x"06ca06c6",	
					x"06c906d1",	x"06dd06de",	x"06aa06e2",	x"06e70717",	
					x"06ee070b",	x"06df06b3",	x"00191031",	x"06bc06a9",	
					x"06c806ab",	x"069706a3",	x"069f06c0",	x"06ac0682",	
					x"06890686",	x"0680069e",	x"067c066b",	x"067f068e",	
					x"06900688",	x"069b06b1",	x"06ae06d2",	x"06d406f0",	
					x"06ef06d2",	x"06d606e9",	x"06cf069c",	x"069f06c4",	
					x"06db06b3",	x"06c406b3",	x"06d006bf",	x"06d406c4",	
					x"06c706b9",	x"06e006da",	x"06d00694",	x"06b206d9",	
					x"06c906d1",	x"06c706b9",	x"06ca06c2",	x"06ee06f2",	
					x"06ea06fc",	x"070306ff",	x"06ee06b3",	x"00192031",	
					x"06b506ab",	x"06aa06af",	x"068806a0",	x"068e069a",	
					x"068c067f",	x"06950696",	x"06980679",	x"06870632",	
					x"06670699",	x"06940697",	x"06ab068f",	x"06b006ad",	
					x"06b706e0",	x"06ee06ec",	x"06b006c0",	x"06b8068e",	
					x"06b006c3",	x"06c906b3",	x"06bc06b3",	x"06bd06d6",	
					x"06cf06cd",	x"06c806d6",	x"06c906ea",	x"06cc069e",	
					x"06c306ca",	x"06a006c8",	x"069e06bf",	x"06d106c4",	
					x"06c906ec",	x"06d80700",	x"06db0712",	x"06e00689",	
					x"00193031",	x"06770688",	x"0673069b",	x"068f06b1",	
					x"068f06a9",	x"067e06bb",	x"06a706b2",	x"068b0668",	
					x"0672065f",	x"065d068f",	x"068006a2",	x"06a106ba",	
					x"06c206f4",	x"06cc06f6",	x"06bd06d5",	x"06d306d9",	
					x"06d8069c",	x"06c506ad",	x"06ad06dd",	x"06d506c1",	
					x"06c306f4",	x"06b606ea",	x"06c606e9",	x"06d006ef",	
					x"06cc06ab",	x"06a906ee",	x"069a06e8",	x"06ab06ec",	
					x"06db0705",	x"06dd0741",	x"06e5071a",	x"06dd0729",	
					x"06f406b5",	x"000a0004",	x"e1380025",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"001a4031",	x"06ac06cd",	x"06a406da",	
					x"06b206ce",	x"06b006d9",	x"06ba06db",	x"069506b4",	
					x"069706a2",	x"06940691",	x"069506dd",	x"06cb06f4",	
					x"06b50702",	x"06d6073e",	x"06d90716",	x"06ea0714",	
					x"07040715",	x"06f206fa",	x"06d30723",	x"07270723",	
					x"07170735",	x"070e072d",	x"0705073b",	x"071b0742",	
					x"07270739",	x"07040720",	x"06fc0736",	x"0710072d",	
					x"070b0722",	x"071c0750",	x"072e078b",	x"07540763",	
					x"07260756",	x"07250707",	x"001a5031",	x"07040713",	
					x"06d50701",	x"06bd070b",	x"06d40717",	x"06c40713",	
					x"06ed072f",	x"06d406f0",	x"06c2070c",	x"06bc0738",	
					x"06fa0745",	x"070f075d",	x"07010757",	x"07120750",	
					x"07460771",	x"07020746",	x"07230722",	x"070b0734",	
					x"07110733",	x"07000741",	x"0716076f",	x"07340775",	
					x"07310763",	x"07210779",	x"0737076c",	x"071c077d",	
					x"073b0775",	x"07120795",	x"072d07a1",	x"072c07e1",	
					x"075c0795",	x"0746077d",	x"073806f6",	x"001a6031",	
					x"06e00712",	x"06de0719",	x"06f70730",	x"06fb0722",	
					x"06e20730",	x"06f3072b",	x"06ca0717",	x"06d106d6",	
					x"06bc0765",	x"07070770",	x"07180774",	x"073a0772",	
					x"074d0764",	x"07680780",	x"0741078f",	x"073d075d",	
					x"0739077d",	x"07410778",	x"076a07a3",	x"075907a4",	
					x"0763079a",	x"07590797",	x"075307a3",	x"07630777",	
					x"075107a6",	x"076c07b2",	x"076207ba",	x"078007f4",	
					x"078307d0",	x"079207d4",	x"079507d1",	x"07790747",	
					x"001a7031",	x"072a074f",	x"07240758",	x"071e0781",	
					x"075a078f",	x"074c077b",	x"073e077a",	x"0731078a",	
					x"0727072f",	x"070507af",	x"077d07b9",	x"076d07ff",	
					x"07920806",	x"07ab07f4",	x"07c107d6",	x"07b60801",	
					x"07a807c2",	x"07ac0800",	x"07b6080d",	x"07ba0810",	
					x"07c40821",	x"07d30819",	x"07f90813",	x"07bb080b",	
					x"07cc07ce",	x"07bc07fd",	x"07f00822",	x"07e50833",	
					x"08110843",	x"08330854",	x"08220851",	x"08290817",	
					x"07f8066b",	x"000a0004",	x"1e285442",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"101b0031",	x"0667067a",	x"067e0682",	
					x"06660659",	x"06610654",	x"064f0638",	x"064d065e",	
					x"0643064d",	x"063205ff",	x"06250632",	x"06640679",	
					x"06810681",	x"068c06a2",	x"06b3068f",	x"06a40683",	
					x"06960677",	x"069d066c",	x"0680066b",	x"066e0659",	
					x"06770664",	x"066c06ba",	x"0674068d",	x"068f0696",	
					x"06a2069d",	x"06a4065d",	x"067d069a",	x"0686069e",	
					x"068606a7",	x"069906a4",	x"068c0699",	x"068d06ab",	
					x"069706d3",	x"06840669",	x"101b1031",	x"0666066d",	
					x"0649066c",	x"064d066c",	x"065e0654",	x"0612064d",	
					x"064a0658",	x"06490616",	x"06620618",	x"0628062d",	
					x"063b0684",	x"067b06a6",	x"06a8068d",	x"068e067f",	
					x"068f06a5",	x"06a3068d",	x"069d0642",	x"06520664",	
					x"06670679",	x"06770686",	x"06af0676",	x"066d068a",	
					x"068d0692",	x"069a0678",	x"068b064f",	x"067d067c",	
					x"06960691",	x"067a0693",	x"06a0068b",	x"0676069e",	
					x"069206a8",	x"06ae06a7",	x"06a0062b",	x"101b2031",	
					x"063d065a",	x"0672066e",	x"06440665",	x"06610654",	
					x"066f0629",	x"063f0645",	x"064a064d",	x"064a061c",	
					x"062f062a",	x"06440640",	x"06480672",	x"066b0687",	
					x"067d0687",	x"0672067b",	x"06870698",	x"06730641",	
					x"0637066b",	x"066c0689",	x"067f0680",	x"0676065e",	
					x"06550679",	x"0676068b",	x"067d067e",	x"06850669",	
					x"06740677",	x"067f068c",	x"068a0675",	x"0676068d",	
					x"066f06aa",	x"0692068a",	x"0673068f",	x"06770637",	
					x"101b3031",	x"0635064f",	x"06410643",	x"0645063b",	
					x"061a063d",	x"06240650",	x"062e0633",	x"06220625",	
					x"061d061f",	x"061f063b",	x"063e064c",	x"065a0671",	
					x"065e067c",	x"06540683",	x"066d0674",	x"066d0687",	
					x"06690650",	x"06360662",	x"06550679",	x"066b0674",	
					x"067e0675",	x"06620683",	x"067b06a1",	x"0690069e",	
					x"06920684",	x"066c0696",	x"0665069d",	x"06710699",	
					x"0695069f",	x"068306aa",	x"068706b2",	x"068606b4",	
					x"0687066e",	x"000a0004",	x"fac7d88a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"101c4031",	x"06490693",	x"065d067a",	
					x"0649066f",	x"06550664",	x"0650067e",	x"06510653",	
					x"06560659",	x"064c065d",	x"063c069a",	x"065f0671",	
					x"066506be",	x"069a06a4",	x"069e06b3",	x"069d06e4",	
					x"06ab0696",	x"0691069b",	x"069606c6",	x"06bb06c6",	
					x"06b306c7",	x"06c106d7",	x"06ca06ce",	x"06b506dd",	
					x"06be06d0",	x"06ad06a1",	x"06a406df",	x"06b406ca",	
					x"06ba06de",	x"06d006ee",	x"06ca06eb",	x"06d306ee",	
					x"06ce06f1",	x"06cf069b",	x"101c5031",	x"069c06a1",	
					x"069006b9",	x"067d06aa",	x"068a06b8",	x"069306ac",	
					x"067c06a9",	x"068f06a5",	x"069706a1",	x"067a06c8",	
					x"06b006d6",	x"06c806d5",	x"06d206f6",	x"06d50701",	
					x"06da06e4",	x"06bb06dd",	x"06bf06d4",	x"06ab0715",	
					x"06ca06e2",	x"06ba06f2",	x"06e006f8",	x"06cb06f5",	
					x"06e10701",	x"06d606fb",	x"06c806e8",	x"06c80725",	
					x"06d50726",	x"06d00729",	x"06f0071d",	x"06ec071e",	
					x"07030723",	x"06fc072b",	x"06f806a3",	x"101c6031",	
					x"06a706d9",	x"069d06d0",	x"06a706ae",	x"069106bb",	
					x"067706cf",	x"06a906c8",	x"068806d2",	x"0684068c",	
					x"068606f7",	x"06c106fe",	x"06e0072f",	x"07120732",	
					x"06c20729",	x"07130721",	x"06f9071b",	x"06f706e3",	
					x"06ee0710",	x"07060718",	x"07000737",	x"070d0738",	
					x"0707073e",	x"07100732",	x"07110732",	x"06e7071a",	
					x"06f20747",	x"07150743",	x"070c0752",	x"0711075a",	
					x"0715075d",	x"07300755",	x"07230741",	x"071606e9",	
					x"101c7031",	x"06d0070a",	x"06f90716",	x"06dc0737",	
					x"07010731",	x"06ed0719",	x"070d0734",	x"06f8070f",	
					x"06da0701",	x"06c10731",	x"071d074e",	x"0732076a",	
					x"077007a5",	x"0758078c",	x"07770799",	x"077a0784",	
					x"07440740",	x"0720077f",	x"075a0781",	x"0761079a",	
					x"077607a0",	x"077107a9",	x"077b07ab",	x"078107b8",	
					x"077e0766",	x"07490799",	x"078307b2",	x"079907c1",	
					x"079207d7",	x"079607cc",	x"07b507da",	x"07ad07ca",	
					x"0799070e",	x"000a0004",	x"344c227f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"201d0031",	x"072f0732",	x"073f071d",	
					x"071206fb",	x"07210719",	x"07170707",	x"06e80717",	
					x"06fa0719",	x"06f90721",	x"07400724",	x"074c0737",	
					x"074d073c",	x"07600748",	x"0768075b",	x"07610760",	
					x"075a0747",	x"0737070c",	x"072d075a",	x"07740754",	
					x"0757073e",	x"0755074d",	x"07420736",	x"0759074f",	
					x"0758075a",	x"075f0732",	x"07510732",	x"072a072f",	
					x"0735074e",	x"0740074e",	x"0744075e",	x"074a0765",	
					x"0729074f",	x"075806f0",	x"201d1031",	x"07320704",	
					x"06d906fe",	x"070906f3",	x"070d0709",	x"06d806e9",	
					x"06ff0703",	x"0705071b",	x"074506cb",	x"06ec0742",	
					x"0742073c",	x"072d075e",	x"07620769",	x"074e074f",	
					x"07600765",	x"076b0731",	x"074506e5",	x"06f30703",	
					x"072c0755",	x"073b072a",	x"07300733",	x"073c0731",	
					x"07440755",	x"0748073f",	x"07520734",	x"073f0743",	
					x"074d0748",	x"0750076b",	x"075c076d",	x"07520761",	
					x"076b0773",	x"07690760",	x"075206f3",	x"201d2031",	
					x"071706fe",	x"07210705",	x"070e0716",	x"06fb06ed",	
					x"06f306e7",	x"06f20712",	x"07010701",	x"071b06e5",	
					x"070006f2",	x"0736074f",	x"075e074d",	x"07530747",	
					x"07510737",	x"07340737",	x"0732074f",	x"073306fc",	
					x"07000749",	x"073b0713",	x"07270739",	x"073a073b",	
					x"073b074e",	x"073e0747",	x"074d0745",	x"07420704",	
					x"07240748",	x"072b0756",	x"072e0733",	x"073a073d",	
					x"07310768",	x"075d0769",	x"07520752",	x"074406dd",	
					x"201d3031",	x"06f406f9",	x"06d70707",	x"06d50718",	
					x"070006f8",	x"06eb06f5",	x"06eb06df",	x"06db070b",	
					x"070206ff",	x"06f70720",	x"070c0741",	x"071f0766",	
					x"07530761",	x"07570756",	x"075a074e",	x"07280743",	
					x"073406f4",	x"070c0733",	x"072f073b",	x"073b075a",	
					x"07620771",	x"073f076e",	x"074f0770",	x"0755074d",	
					x"073e0754",	x"073c0784",	x"074b075c",	x"072b076b",	
					x"07280764",	x"07390786",	x"074e0793",	x"075c0796",	
					x"07580724",	x"000a0004",	x"9d4d3a02",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"201e4031",	x"071a0730",	x"0742072e",	
					x"071b072e",	x"072d0745",	x"0701070a",	x"0724073c",	
					x"07000741",	x"0720072c",	x"0729074f",	x"07610772",	
					x"07680776",	x"076907a3",	x"075b0790",	x"07660783",	
					x"07810773",	x"0764075a",	x"07520796",	x"07690799",	
					x"078407ad",	x"0791079a",	x"077c07c4",	x"079607c4",	
					x"07aa07c2",	x"079f0798",	x"079907c0",	x"07b807a6",	
					x"079e07b9",	x"078c07a3",	x"078207c2",	x"079c07cf",	
					x"07af07c8",	x"07920747",	x"201e5031",	x"0744076a",	
					x"0748079d",	x"074b078b",	x"0745076a",	x"0732076c",	
					x"074e0788",	x"0756077b",	x"07550792",	x"078307c9",	
					x"078607d3",	x"079107b7",	x"07a707ba",	x"07ad07d7",	
					x"07b607b1",	x"07ac07bf",	x"07850790",	x"076307db",	
					x"079807e0",	x"078b07e1",	x"07a007f4",	x"079507dc",	
					x"07c20802",	x"07a507e8",	x"07b007cc",	x"07ab07f9",	
					x"07c007e4",	x"07aa07ea",	x"07950803",	x"07aa0806",	
					x"07be080d",	x"07c407e3",	x"07a40765",	x"201e6031",	
					x"077107a7",	x"07850789",	x"0760077a",	x"075307a7",	
					x"075c0774",	x"074407c7",	x"076d079e",	x"077b07ae",	
					x"077907fc",	x"07bf0802",	x"07b207f1",	x"07bf0807",	
					x"07be080a",	x"07eb0800",	x"07d907e5",	x"07d907e7",	
					x"07c607f4",	x"07e6080a",	x"07d7081b",	x"07f1082a",	
					x"07df0823",	x"07f30833",	x"07e2082f",	x"07e60801",	
					x"07f30821",	x"07db082b",	x"07ce0852",	x"07e6083b",	
					x"07fc0841",	x"07fd0842",	x"07fc0838",	x"07e807c9",	
					x"201e7031",	x"07b507f7",	x"07b107d2",	x"079d07ef",	
					x"07ac0810",	x"07a007f5",	x"0794081b",	x"079c0816",	
					x"07b507f3",	x"07d7085f",	x"0829086d",	x"08270870",	
					x"0824087c",	x"082e088a",	x"0856086c",	x"0843086a",	
					x"0845087a",	x"082c0886",	x"084608a8",	x"085b08a0",	
					x"085808a2",	x"084908a3",	x"08670887",	x"085408d7",	
					x"086f0881",	x"087c08a9",	x"087f0896",	x"087308b9",	
					x"088808b8",	x"088708bf",	x"088708d2",	x"0895088e",	
					x"089f06ff",	x"000a0004",	x"dfbc92bd",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"301f0031",	x"06f006e6",	x"06df0709",	
					x"06fb06ea",	x"072706ef",	x"06fa070a",	x"06f106fa",	
					x"06e206f3",	x"06ef06c8",	x"06d906ff",	x"07230730",	
					x"072a0711",	x"07210755",	x"073a075e",	x"0751075b",	
					x"07430711",	x"071106de",	x"070a0711",	x"0727071d",	
					x"071606ee",	x"071b0744",	x"07320748",	x"07420749",	
					x"0715071d",	x"070f0718",	x"071f071b",	x"0724071c",	
					x"070c070f",	x"070f070c",	x"0701072f",	x"072d074f",	
					x"0749073a",	x"071306d0",	x"301f1031",	x"06f006c6",	
					x"06e506cc",	x"06c506cf",	x"06bc06d1",	x"06bd06d1",	
					x"06ef06d6",	x"06c506dd",	x"06df06b1",	x"06c80714",	
					x"071b073b",	x"07480723",	x"07370719",	x"071c0711",	
					x"071b071c",	x"07150719",	x"071406c5",	x"06db071c",	
					x"07210709",	x"07150727",	x"07360739",	x"07480720",	
					x"073f0754",	x"0740072c",	x"072f0713",	x"070c070d",	
					x"070d0739",	x"0743072f",	x"07250712",	x"07070722",	
					x"07180724",	x"07210725",	x"073e06dc",	x"301f2031",	
					x"06e306d3",	x"06d306b7",	x"06ba06bd",	x"06cc06d6",	
					x"06e906cd",	x"06c506d5",	x"06ce06e4",	x"07090677",	
					x"06e10709",	x"0723070f",	x"071e071e",	x"07090710",	
					x"071f0728",	x"07230723",	x"0703070b",	x"070e06db",	
					x"07080709",	x"0705070a",	x"06fd0703",	x"0718071f",	
					x"0719072b",	x"07250746",	x"0736072c",	x"072006e6",	
					x"06f1070f",	x"07210739",	x"07080712",	x"07050731",	
					x"07100708",	x"0703071f",	x"0709072e",	x"0722069f",	
					x"301f3031",	x"069606b0",	x"06a806e5",	x"06be06ba",	
					x"06c0070c",	x"06c506e2",	x"06cf06d5",	x"06cd06d5",	
					x"06c806de",	x"06d606f3",	x"06fd0703",	x"06f70727",	
					x"07100724",	x"0705071f",	x"070d06eb",	x"06ea06f6",	
					x"070a06de",	x"06db06f9",	x"06f106ff",	x"06f3072c",	
					x"07270733",	x"071e0726",	x"0728075a",	x"07080753",	
					x"07240729",	x"07100732",	x"07170718",	x"0702071a",	
					x"0700072d",	x"0702072f",	x"07020739",	x"06eb072f",	
					x"070d06e1",	x"000a0004",	x"c758246f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"30204031",	x"06b206f7",	x"06f206ee",	
					x"06cd06f0",	x"06ca0706",	x"06d906f4",	x"06ee0700",	
					x"070e070f",	x"07090707",	x"06f80731",	x"0736073f",	
					x"0733074c",	x"07420751",	x"073d0752",	x"0735075b",	
					x"0739072c",	x"07170708",	x"06f90759",	x"07400754",	
					x"073c0757",	x"0752077c",	x"07490769",	x"074d0771",	
					x"075c0774",	x"07570743",	x"0744074f",	x"073b077f",	
					x"0759075e",	x"0765076f",	x"07510779",	x"075c0783",	
					x"074e0776",	x"07440748",	x"30205031",	x"0722074b",	
					x"0727073b",	x"06f70748",	x"072b074c",	x"0720074f",	
					x"072c076a",	x"0750076f",	x"0751075b",	x"0756077e",	
					x"0788077a",	x"076a077b",	x"07660776",	x"0759078b",	
					x"0773077e",	x"07750775",	x"075b0750",	x"072507a8",	
					x"074d078d",	x"0769079b",	x"077f07bd",	x"077307b0",	
					x"077507c1",	x"077d07c8",	x"077a07a4",	x"075907e1",	
					x"078507a6",	x"077907b0",	x"078107a3",	x"074707d4",	
					x"077b07d0",	x"079307c1",	x"07910738",	x"30206031",	
					x"070b0766",	x"073c0763",	x"072e0762",	x"07440757",	
					x"074f075d",	x"0759075e",	x"07400757",	x"074e0772",	
					x"075607bd",	x"079e07c2",	x"079907bd",	x"07b307c7",	
					x"07a307b3",	x"077707b8",	x"078507c7",	x"07890790",	
					x"078507bc",	x"078c07e7",	x"078f07ec",	x"07b707ec",	
					x"07b007fd",	x"07a50801",	x"07a807e4",	x"07a807c0",	
					x"07af07f2",	x"07d207dc",	x"07ad07e6",	x"07c10814",	
					x"07ad07ff",	x"07e00813",	x"07c70800",	x"07c8078a",	
					x"30207031",	x"076f0797",	x"074c07a8",	x"076007b1",	
					x"078007f5",	x"078f07b8",	x"077d07d4",	x"079407e1",	
					x"07d307f1",	x"07cd084a",	x"07e00842",	x"0806082d",	
					x"08000823",	x"07f6084b",	x"0827083b",	x"0807081c",	
					x"07f607e4",	x"07e6083b",	x"08180858",	x"08030862",	
					x"0839085c",	x"08180868",	x"083d0886",	x"085d0872",	
					x"0848082d",	x"082a086d",	x"085b087d",	x"081d086a",	
					x"084e08ba",	x"0854089e",	x"086a088c",	x"086d086d",	
					x"085206c8",	x"000a0004",	x"05ed754a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0121002e",	x"06650669",	x"065c0655",	
					x"065b0663",	x"065e0653",	x"064b0663",	x"0636065b",	
					x"0662065c",	x"0659065d",	x"0659065e",	x"0675069e",	
					x"06830662",	x"067d0662",	x"06580672",	x"0686069d",	
					x"067e068f",	x"068a063e",	x"06540669",	x"06980678",	
					x"0675069c",	x"067d067f",	x"067c0665",	x"067b06a5",	
					x"068d066a",	x"066f064b",	x"065e0672",	x"067b06a6",	
					x"068c0696",	x"06a106a4",	x"0694067c",	x"068206c2",	
					x"068d0683",	x"06750671",	x"0121102e",	x"0666063c",	
					x"0655063e",	x"06320640",	x"064e0617",	x"06220620",	
					x"062a0634",	x"0630063d",	x"065b0623",	x"06500656",	
					x"0668066c",	x"0663066e",	x"066d0674",	x"068a0663",	
					x"067f0678",	x"06830678",	x"066a0632",	x"064f0673",	
					x"067d0664",	x"065b064a",	x"06690678",	x"0683067f",	
					x"0685067b",	x"066d0670",	x"06700632",	x"06650660",	
					x"068b066e",	x"0684068a",	x"0692068a",	x"067e068a",	
					x"06b8068d",	x"06990681",	x"06810626",	x"0121202e",	
					x"06230629",	x"063c062a",	x"063c0612",	x"06430623",	
					x"063a0629",	x"064b0652",	x"0657065d",	x"0663061f",	
					x"063b0633",	x"06540638",	x"06470660",	x"0651064f",	
					x"066e0674",	x"068a0682",	x"067c0678",	x"06860641",	
					x"06510639",	x"065a0635",	x"063d0654",	x"066a0654",	
					x"064f0670",	x"0662066f",	x"065b0661",	x"064f063a",	
					x"06560658",	x"064e0645",	x"06510670",	x"066e068f",	
					x"067d065f",	x"0673068c",	x"066a0679",	x"06600615",	
					x"0121302e",	x"060f0628",	x"0623061d",	x"0621061d",	
					x"060f0602",	x"06010627",	x"06300639",	x"0636062b",	
					x"0634061a",	x"063b064c",	x"06620660",	x"064a065c",	
					x"06610649",	x"063a0644",	x"06530667",	x"0651064a",	
					x"06540621",	x"063a063f",	x"0651064e",	x"06420643",	
					x"06650669",	x"06610681",	x"06770661",	x"065e0677",	
					x"06520643",	x"064e0666",	x"06590687",	x"065d0676",	
					x"06720672",	x"06680686",	x"066c0687",	x"065b0675",	
					x"06610626",	x"000a0004",	x"b865cd8c",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0122402e",	x"0613063a",	x"06360653",	
					x"0619061a",	x"062a062e",	x"063c0638",	x"063b0661",	
					x"06540656",	x"06420654",	x"06590654",	x"065a067b",	
					x"0651065e",	x"06760666",	x"0668067a",	x"0663066f",	
					x"06800677",	x"067b0652",	x"065d066f",	x"06770682",	
					x"067b068f",	x"0699068c",	x"06890696",	x"06a4069b",	
					x"0689065f",	x"0680067c",	x"068c067a",	x"068906a2",	
					x"06a306a7",	x"06c1069d",	x"069106ad",	x"06a606ba",	
					x"06a306a4",	x"069b066e",	x"0122502e",	x"06590689",	
					x"06730655",	x"0647064f",	x"0640066e",	x"06410676",	
					x"06680668",	x"06670694",	x"0681066b",	x"0682069a",	
					x"068c069f",	x"06910693",	x"069c06ac",	x"06a1069b",	
					x"06a7069b",	x"069906a3",	x"06920680",	x"066b0688",	
					x"069a06af",	x"068f06a2",	x"069d06ab",	x"06b206b5",	
					x"068f06ad",	x"06a706b1",	x"06a306a3",	x"069606ca",	
					x"06b306d5",	x"06bd06e2",	x"06ad06e4",	x"06b906d5",	
					x"06b006da",	x"06bc06c8",	x"06b10671",	x"0122602e",	
					x"065b0686",	x"066c0689",	x"06730653",	x"06630667",	
					x"066b06a2",	x"06ab067b",	x"0668067d",	x"068f067a",	
					x"066f068f",	x"067e06c4",	x"06a2069e",	x"06a506cf",	
					x"06d206d2",	x"06cc06fc",	x"06cb06c9",	x"06d306b2",	
					x"06a606c7",	x"06c106d4",	x"06b306df",	x"06d906e2",	
					x"06dd06ec",	x"06e006e4",	x"06d306f1",	x"06c606c7",	
					x"06d60709",	x"07000700",	x"06e60709",	x"06f30702",	
					x"06db070a",	x"06f40713",	x"06eb0702",	x"06ec069c",	
					x"0122702e",	x"065a0696",	x"06880699",	x"0673068e",	
					x"067806a1",	x"067d06b4",	x"069e06c2",	x"06c80694",	
					x"068606c2",	x"06a306c2",	x"0706071c",	x"06f806f9",	
					x"06d6071a",	x"06f9073b",	x"07140741",	x"06fa0723",	
					x"071f06e7",	x"06ea074b",	x"071c0722",	x"0724073c",	
					x"07370754",	x"07470757",	x"0746073e",	x"072d0743",	
					x"07300729",	x"0738074e",	x"074b076a",	x"075c074a",	
					x"075a0777",	x"07640776",	x"075b0780",	x"07560769",	
					x"0754071b",	x"000a0004",	x"deabfcdd",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1123002e",	x"07110729",	x"07100733",	
					x"07250700",	x"071b06fa",	x"07120728",	x"0720076a",	
					x"074d0762",	x"07500726",	x"0728075f",	x"07720789",	
					x"0776077a",	x"077a076e",	x"07500734",	x"07500745",	
					x"0750074b",	x"0774072f",	x"074f0748",	x"0755075e",	
					x"07550742",	x"074c0742",	x"07470740",	x"074d075e",	
					x"075b0750",	x"0748070d",	x"076b0767",	x"0772075e",	
					x"075c0762",	x"07670769",	x"075e0750",	x"07710787",	
					x"074c075d",	x"074106ec",	x"1123102e",	x"06e606f8",	
					x"073b0722",	x"07260715",	x"071a0704",	x"070d0700",	
					x"06fe0710",	x"0719073b",	x"07430713",	x"07230749",	
					x"074c074e",	x"073e0752",	x"07440737",	x"0739072c",	
					x"073e074c",	x"0743073a",	x"073a0726",	x"07280742",	
					x"076d0750",	x"07430758",	x"0750071e",	x"07350722",	
					x"071f073f",	x"07380756",	x"0767071f",	x"07490753",	
					x"075a0768",	x"07520762",	x"075a0742",	x"075d0737",	
					x"074d0744",	x"07400758",	x"0748070c",	x"1123202e",	
					x"06f306fb",	x"06f80702",	x"070606d4",	x"06ee0718",	
					x"071d06fb",	x"072606e9",	x"070e06f7",	x"072406e4",	
					x"070a0732",	x"075a072c",	x"07430726",	x"072e0719",	
					x"072b0718",	x"072f0715",	x"0725071d",	x"073b06f9",	
					x"0713072d",	x"072b0724",	x"0727071d",	x"07280707",	
					x"070b0724",	x"071f071f",	x"071b0730",	x"073f071a",	
					x"07360734",	x"072f0735",	x"073b072d",	x"07390736",	
					x"07260734",	x"072d0731",	x"072b0725",	x"071006c6",	
					x"1123302e",	x"06b806cf",	x"06b706e4",	x"06d206d5",	
					x"06c906ec",	x"06ed06e1",	x"06ef06b8",	x"06ca0719",	
					x"070706e6",	x"06f4071e",	x"0719071c",	x"070d072b",	
					x"070d06f3",	x"07180727",	x"071f0730",	x"07310722",	
					x"071106fb",	x"06ff0729",	x"07130727",	x"07180721",	
					x"0718071d",	x"0719071d",	x"07020731",	x"0713074c",	
					x"072a06fa",	x"07320728",	x"07330743",	x"07190739",	
					x"072b073f",	x"07340753",	x"0730075c",	x"07230755",	
					x"072f06e8",	x"000a0004",	x"5f0534b0",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1124402e",	x"06d306f8",	x"06ec0702",	
					x"06ef06ed",	x"06fc0706",	x"06ed0704",	x"07020700",	
					x"07150710",	x"071c0704",	x"071d0716",	x"071a0737",	
					x"073e0740",	x"07320745",	x"073e073a",	x"073e0742",	
					x"0749074b",	x"0750073d",	x"07510753",	x"07800754",	
					x"0747077f",	x"0766075d",	x"076c075b",	x"07510753",	
					x"0760074f",	x"07480751",	x"075d076b",	x"0761078b",	
					x"0771077a",	x"076b078c",	x"0775078e",	x"077607a6",	
					x"07760771",	x"074f073d",	x"1124502e",	x"071c072b",	
					x"07000742",	x"07110750",	x"07090747",	x"07210747",	
					x"073b073e",	x"072b074c",	x"074b074f",	x"074c077b",	
					x"07600783",	x"0750076b",	x"07650771",	x"0774077a",	
					x"076d076d",	x"0764077e",	x"076f0769",	x"075c077b",	
					x"077e078c",	x"076b077a",	x"07630785",	x"076a079e",	
					x"077d07a7",	x"077807a3",	x"077d0794",	x"077a07b8",	
					x"078a07ae",	x"078107bd",	x"078e07c3",	x"078c07b6",	
					x"078c07d3",	x"079e07ad",	x"077e073c",	x"1124602e",	
					x"0719072e",	x"06fa074d",	x"07280756",	x"0732075f",	
					x"07350747",	x"070a0760",	x"0748075b",	x"07430774",	
					x"0764077c",	x"0756078f",	x"077007b4",	x"077f07b4",	
					x"077507ab",	x"077b0793",	x"077a0794",	x"0784079e",	
					x"078d079e",	x"07a807b8",	x"07a007b6",	x"07c307af",	
					x"07c007bf",	x"07ac07cc",	x"07a907ac",	x"079f07c6",	
					x"07bd07eb",	x"07dd07e4",	x"07bc07bc",	x"07a407f1",	
					x"07cd07f7",	x"07c107e4",	x"07bd07e2",	x"0791076d",	
					x"1124702e",	x"0761078b",	x"0768077b",	x"0744078f",	
					x"07700789",	x"07430780",	x"076d07af",	x"07a9079e",	
					x"079707ab",	x"079607b7",	x"07b407ea",	x"07c407f1",	
					x"07e60803",	x"07cb07f1",	x"07f3080d",	x"07e907ed",	
					x"07ec07e8",	x"07e607f9",	x"07eb07ef",	x"07e6083e",	
					x"07f40848",	x"07fd0821",	x"080e081d",	x"081a082c",	
					x"083507e9",	x"08000864",	x"08260869",	x"0830083f",	
					x"08430867",	x"082c0891",	x"08370851",	x"08440842",	
					x"082106ed",	x"000a0004",	x"876569ee",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2125002e",	x"06db06c9",	x"06bf06b3",	
					x"06a60694",	x"06a506b6",	x"06c406d4",	x"06e106fa",	
					x"072806d8",	x"06e806e1",	x"06d606f7",	x"06fd0710",	
					x"06eb070c",	x"07280717",	x"07140706",	x"06ff06f0",	
					x"06fa06f8",	x"06f806d7",	x"070d06f1",	x"070b06ee",	
					x"070206f5",	x"071506f3",	x"06f406f1",	x"070006f9",	
					x"06ff06fa",	x"06ec06f5",	x"06f20722",	x"07150705",	
					x"0700071e",	x"06f8072c",	x"070f0708",	x"06f506fc",	
					x"06e60701",	x"06f106a4",	x"2125102e",	x"069d0690",	
					x"068c06b9",	x"06c006a3",	x"06a50692",	x"068306b2",	
					x"06ce06d5",	x"06be06e1",	x"06b306b4",	x"06d306e6",	
					x"06e106ec",	x"06ed06df",	x"06d306de",	x"06de06d9",	
					x"06e006d9",	x"06eb06ce",	x"06f406c1",	x"06c506e8",	
					x"06e506df",	x"06f106e3",	x"070606e5",	x"06fa06ee",	
					x"071706eb",	x"06d506ed",	x"06fe06e2",	x"06fc070c",	
					x"07380707",	x"07010709",	x"071706dc",	x"06e10715",	
					x"07040712",	x"070d06f8",	x"06e506a8",	x"2125202e",	
					x"069e0691",	x"069506a6",	x"06a30681",	x"06a106ae",	
					x"06d106a4",	x"06be06aa",	x"069c06a0",	x"06b30689",	
					x"069a06c1",	x"06ea06c0",	x"06ce06d9",	x"06ef06d8",	
					x"06d606d6",	x"06da06df",	x"06e006e2",	x"06c606ac",	
					x"06bd06ca",	x"06dd06ea",	x"06c706de",	x"06ef06da",	
					x"06cd06db",	x"06da06e6",	x"06e906dd",	x"06c506c6",	
					x"06cd06e4",	x"06de06f8",	x"06e906ee",	x"06f506fc",	
					x"06ce06e5",	x"06cf06e3",	x"06cd06c5",	x"06cc0662",	
					x"2125302e",	x"06860675",	x"06670680",	x"066a068f",	
					x"069506ac",	x"068f06ae",	x"0699069a",	x"06a406aa",	
					x"06a80693",	x"069606c5",	x"06bf06e9",	x"06e706c4",	
					x"06c106cf",	x"06b306c7",	x"06d406cd",	x"06c906cc",	
					x"06c00692",	x"06a706cf",	x"06d806dc",	x"06e206d2",	
					x"06e306c5",	x"06c506ce",	x"06d306e1",	x"06d406e7",	
					x"06c006bb",	x"06db06f5",	x"06de06f4",	x"06e606e8",	
					x"06e10704",	x"06e506ef",	x"06de06f6",	x"06d906f0",	
					x"06d3067d",	x"000a0004",	x"74150a63",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2126402e",	x"066d0688",	x"06a906bb",	
					x"06b206a5",	x"06a506ab",	x"06b306ca",	x"06ab06c2",	
					x"06a606e0",	x"06d1069e",	x"06ae06df",	x"06ca06e6",	
					x"070106cb",	x"06e80715",	x"070b06fc",	x"06fa06fe",	
					x"070706e7",	x"06f106d1",	x"06da06f7",	x"071d071a",	
					x"071a0704",	x"070706fe",	x"072e0707",	x"070106f9",	
					x"07010705",	x"06fc06fc",	x"0704071a",	x"0725071d",	
					x"07090734",	x"07320724",	x"07200726",	x"07280730",	
					x"071f072b",	x"071906a9",	x"2126502e",	x"06af06d8",	
					x"06c706df",	x"06d906da",	x"06cb06f7",	x"06eb0701",	
					x"06e906f9",	x"06f70708",	x"070706e8",	x"06ea0701",	
					x"06f7072e",	x"070f0715",	x"073f071e",	x"0717070f",	
					x"0718071a",	x"06fe0715",	x"070306f9",	x"06f20717",	
					x"0730071b",	x"070f071f",	x"0712073b",	x"0702073d",	
					x"071c0743",	x"07250742",	x"0739073e",	x"07290747",	
					x"07320740",	x"072c0750",	x"072e0755",	x"073a0749",	
					x"073f0759",	x"072d076b",	x"073a06d2",	x"2126602e",	
					x"06a006d4",	x"06d6071c",	x"06f506f0",	x"06f006f0",	
					x"06d606f5",	x"06f6071d",	x"06fc06f6",	x"06f306d8",	
					x"06f9072d",	x"0723072d",	x"07290736",	x"07290739",	
					x"07220762",	x"074d0755",	x"07420739",	x"07230725",	
					x"071c074e",	x"07520768",	x"0742072d",	x"073d0763",	
					x"07540762",	x"075a0774",	x"07480766",	x"07370759",	
					x"07490789",	x"075f0790",	x"07610778",	x"075e0796",	
					x"0756079c",	x"07750794",	x"075c0791",	x"0749072c",	
					x"2126702e",	x"06ef0705",	x"06c00714",	x"06f60724",	
					x"0722076f",	x"0718070a",	x"07060731",	x"07200763",	
					x"071a0758",	x"07520778",	x"07640791",	x"077c0790",	
					x"079f07a2",	x"076c0790",	x"078c07e1",	x"0778078e",	
					x"076c0772",	x"07790796",	x"07b207bd",	x"07ab07c4",	
					x"07ba07eb",	x"07b707c4",	x"07a907c1",	x"07a107d0",	
					x"07a307d6",	x"07bf07ec",	x"07e207e9",	x"07ea07f4",	
					x"07f10817",	x"07eb0819",	x"07e60817",	x"07dc0808",	
					x"07ca06de",	x"000a0004",	x"9d2b3ce5",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3127002e",	x"06e7070c",	x"0717070b",	
					x"070a06ef",	x"06ef070b",	x"07130707",	x"070e070d",	
					x"071d0718",	x"07210700",	x"0729072d",	x"072c0729",	
					x"0730072a",	x"0777075f",	x"073f075e",	x"07510730",	
					x"073c0719",	x"070c06f8",	x"06f80722",	x"073a0758",	
					x"07540753",	x"0759073d",	x"072f0741",	x"0750075f",	
					x"0770073b",	x"071606d4",	x"0710072c",	x"07400750",	
					x"0730074f",	x"07610777",	x"07640752",	x"07440760",	
					x"0726072b",	x"072106d7",	x"3127102e",	x"06e706dd",	
					x"06f606dc",	x"06e106cb",	x"06f706e9",	x"06f006d2",	
					x"07010701",	x"07120716",	x"070406d3",	x"0713074c",	
					x"073b0742",	x"0749073b",	x"0759074b",	x"074e072d",	
					x"075b0736",	x"07370717",	x"072306c3",	x"06e30717",	
					x"07400709",	x"072d0735",	x"0754072b",	x"0729071f",	
					x"072d0714",	x"07210727",	x"0732071a",	x"072c0730",	
					x"072e0732",	x"0747072f",	x"07400750",	x"07450745",	
					x"07390740",	x"0740072b",	x"073306eb",	x"3127202e",	
					x"06e506c4",	x"06fd06c4",	x"06ff06c0",	x"06d906e6",	
					x"06f506d3",	x"06fc06f9",	x"071706b4",	x"070806a9",	
					x"06d20710",	x"07360710",	x"07290703",	x"07130712",	
					x"071c0715",	x"07290724",	x"06ef06fe",	x"070c06b6",	
					x"0707070a",	x"0721070d",	x"071a0715",	x"06f70719",	
					x"070c071a",	x"071a0738",	x"0712071f",	x"06f206be",	
					x"06e5071c",	x"072b071e",	x"07390715",	x"07270713",	
					x"07220748",	x"07280742",	x"0707070e",	x"06df06bf",	
					x"3127302e",	x"06ac06d3",	x"06ba06e5",	x"06cf06cc",	
					x"06c506bd",	x"06c806da",	x"06c306df",	x"06c606e3",	
					x"06e706e3",	x"06d106d9",	x"06dc070e",	x"06f60708",	
					x"06ef0710",	x"06fe0705",	x"06fa070c",	x"06fd0709",	
					x"070406ce",	x"06e506f0",	x"07060705",	x"0712071a",	
					x"071c0708",	x"0721071f",	x"070d071c",	x"070a06fe",	
					x"0702070a",	x"070e0702",	x"07250720",	x"07080725",	
					x"07060722",	x"07260734",	x"071e073d",	x"07190729",	
					x"070e06bc",	x"000a0004",	x"d344274e",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3128402e",	x"06b706d4",	x"06bc06d1",	
					x"06ca06cf",	x"06d206d6",	x"06c60700",	x"06e00704",	
					x"070806ff",	x"0711070a",	x"06fc0718",	x"07290727",	
					x"071a0726",	x"07370739",	x"070f072d",	x"072d0726",	
					x"07180712",	x"06f1072a",	x"0706072c",	x"07320730",	
					x"072d0733",	x"07560759",	x"07460748",	x"0751073c",	
					x"07290734",	x"072b0734",	x"073d0740",	x"0745075f",	
					x"0754075e",	x"0779078a",	x"0758075d",	x"075d0756",	
					x"07430763",	x"07560708",	x"3128502e",	x"06d10701",	
					x"07000713",	x"07030716",	x"070d06ff",	x"07070734",	
					x"07230753",	x"0764075a",	x"07530705",	x"07260755",	
					x"07560758",	x"074f0760",	x"076c0767",	x"07440775",	
					x"0764074d",	x"074f0739",	x"0734071f",	x"07260772",	
					x"0763077b",	x"07540770",	x"077a078a",	x"076c0767",	
					x"0765077e",	x"07600766",	x"07320760",	x"075007b6",	
					x"077307af",	x"076a07b1",	x"077807b8",	x"078f078f",	
					x"076307b4",	x"0775076e",	x"07320722",	x"3128602e",	
					x"07050745",	x"06df0737",	x"07300736",	x"07140738",	
					x"070c0766",	x"074f074a",	x"07380740",	x"072d072d",	
					x"07220783",	x"077c0783",	x"076c078f",	x"07720794",	
					x"077c0790",	x"07540797",	x"07620787",	x"07600785",	
					x"07600786",	x"07880791",	x"07790796",	x"078707c0",	
					x"077c079d",	x"079007c0",	x"079207ab",	x"07a00788",	
					x"078b07e7",	x"07be07e8",	x"07b507dd",	x"07bb07cf",	
					x"079d07d9",	x"078907c3",	x"077d07c5",	x"0781074d",	
					x"3128702e",	x"0755075c",	x"07480772",	x"07560755",	
					x"074b0788",	x"07330787",	x"073d07b3",	x"079e078c",	
					x"0777078d",	x"078507ca",	x"07ad080d",	x"07ce07ca",	
					x"07b007f5",	x"07b207e6",	x"07e107e4",	x"07dc07c9",	
					x"07ae07ec",	x"07db07f5",	x"08010808",	x"07fa07fd",	
					x"07fa0844",	x"07e10813",	x"080b080a",	x"07da07fe",	
					x"07f6080e",	x"080e080c",	x"080e0834",	x"08260828",	
					x"08220868",	x"08140856",	x"08380844",	x"07fe082f",	
					x"0800065e",	x"000a0004",	x"fb3b5d5b",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0129002f",	x"0668067b",	x"06780686",	
					x"067a0667",	x"0643066c",	x"065a0656",	x"063f0644",	
					x"062e0641",	x"06610644",	x"06540660",	x"06650685",	
					x"066e069f",	x"06ad0695",	x"068c0689",	x"068e0691",	
					x"06950688",	x"069c063d",	x"06700688",	x"06850683",	
					x"06830697",	x"069d068b",	x"067f0691",	x"06950693",	
					x"069a0699",	x"0692063c",	x"06780692",	x"06b10695",	
					x"06b206a5",	x"06ad068a",	x"066e0694",	x"069c06aa",	
					x"06ac06a8",	x"06950667",	x"0129102f",	x"06540626",	
					x"06460661",	x"063d0651",	x"06400633",	x"063a0637",	
					x"0623063a",	x"0626063d",	x"063a0620",	x"064e0653",	
					x"0666068e",	x"068a0688",	x"0678066a",	x"068f0689",	
					x"06900682",	x"06730669",	x"066e064a",	x"064d0684",	
					x"067d0675",	x"067d0678",	x"06960696",	x"06a6068d",	
					x"0685067a",	x"068b068c",	x"0696063a",	x"067e067a",	
					x"068b0688",	x"069a0689",	x"0688067b",	x"0668068b",	
					x"06a2069f",	x"06a4068d",	x"06ac063e",	x"0129202f",	
					x"062f0642",	x"0640066a",	x"0659064a",	x"064f0659",	
					x"06550620",	x"061e062d",	x"0631061e",	x"064205f4",	
					x"063f0658",	x"067b0657",	x"06650666",	x"0671066a",	
					x"066e0665",	x"067c0671",	x"06730689",	x"066c063a",	
					x"06540665",	x"06600676",	x"0668067a",	x"06a1065a",	
					x"0667066d",	x"065b065b",	x"065e0662",	x"0661065d",	
					x"066e0675",	x"0667066e",	x"0668066f",	x"0678068f",	
					x"067f0679",	x"06800698",	x"06780697",	x"06860615",	
					x"0129302f",	x"06230627",	x"06210635",	x"062c063f",	
					x"0630062b",	x"0609061c",	x"06130616",	x"06040611",	
					x"06220625",	x"0625065e",	x"06320662",	x"063a0663",	
					x"06750671",	x"065b0651",	x"0658064f",	x"064b0675",	
					x"064f0655",	x"06540660",	x"0656066b",	x"064f0666",	
					x"06790669",	x"064b068a",	x"06750684",	x"0670068b",	
					x"0666065c",	x"064f066a",	x"0662069a",	x"066a069e",	
					x"067c0693",	x"0679069e",	x"067906a2",	x"0698069e",	
					x"06850654",	x"000a0004",	x"bcffd441",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"012a402f",	x"06400644",	x"0646064b",	
					x"063f0648",	x"0625063d",	x"060b0639",	x"0657064e",	
					x"061b064b",	x"0630064a",	x"06540681",	x"068d0686",	
					x"06660686",	x"068d0673",	x"06540684",	x"068c068b",	
					x"067b068d",	x"066b0689",	x"067606b2",	x"06bf06bd",	
					x"06c106b3",	x"06af06c9",	x"06a806cd",	x"06a406b4",	
					x"06a906aa",	x"06a70695",	x"069406cb",	x"06a806cf",	
					x"06aa06dd",	x"06d606ca",	x"069c06cf",	x"06bf06dd",	
					x"06be06c3",	x"06b00669",	x"012a502f",	x"066c0684",	
					x"068a067d",	x"06830689",	x"066f068f",	x"06630683",	
					x"0669067c",	x"06820685",	x"066b067c",	x"065f06b5",	
					x"06c106c1",	x"06b906ba",	x"06a006cd",	x"06b706c1",	
					x"06b606cf",	x"06b706d9",	x"06a006bc",	x"06a006d0",	
					x"06b306d0",	x"06af06c6",	x"06b906f5",	x"06be06e2",	
					x"06b206eb",	x"06d506e5",	x"06c406c9",	x"06b9070b",	
					x"06c8070c",	x"06eb070c",	x"06d3070f",	x"06e1070c",	
					x"06dc071e",	x"06e706dd",	x"06c6067e",	x"012a602f",	
					x"0646068b",	x"065a06ad",	x"06970690",	x"067e067b",	
					x"065f06ae",	x"067e06a1",	x"065f068c",	x"0667069a",	
					x"067906d3",	x"069f06c3",	x"06ac06df",	x"06da06db",	
					x"06e20708",	x"06ec0702",	x"06c706ef",	x"06e606f1",	
					x"06e306ef",	x"06e806f5",	x"06d40704",	x"06f50720",	
					x"06e0071d",	x"06f30731",	x"06f20738",	x"06fc06fd",	
					x"06e90711",	x"06ed0719",	x"06e60727",	x"06f10726",	
					x"0703074e",	x"0706074e",	x"07090729",	x"06f5068e",	
					x"012a702f",	x"066006b5",	x"06860703",	x"06b306a3",	
					x"069206c8",	x"068606fb",	x"069306fd",	x"069706ea",	
					x"06a406af",	x"06830715",	x"06e90769",	x"071b072f",	
					x"06f6075a",	x"06f0073a",	x"0713074a",	x"071b076c",	
					x"07250722",	x"071b0760",	x"07270757",	x"0727076a",	
					x"072e07a4",	x"07220760",	x"074b0748",	x"072b0760",	
					x"072f0748",	x"073e0770",	x"074c078a",	x"0748078b",	
					x"077107cd",	x"0794079c",	x"078e07b6",	x"07770779",	
					x"0756075a",	x"000a0004",	x"e7231019",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"112b002f",	x"0756077a",	x"07670792",	
					x"0772075e",	x"076f075c",	x"074c074b",	x"07590741",	
					x"07250713",	x"06f406ee",	x"06f306fb",	x"06f2071f",	
					x"0725074e",	x"074a074c",	x"075a0765",	x"077a0782",	
					x"07840755",	x"076f0740",	x"0739074a",	x"0751075a",	
					x"07570760",	x"07690761",	x"07570768",	x"07820759",	
					x"075f0763",	x"0785072e",	x"0747074c",	x"075a074e",	
					x"07540766",	x"0778078f",	x"0742075e",	x"075a0776",	
					x"0765077d",	x"07590738",	x"112b102f",	x"0733072f",	
					x"073d0774",	x"075f0752",	x"073c074b",	x"072d0751",	
					x"073806fc",	x"07040703",	x"06fc06ef",	x"06e206d3",	
					x"06e70707",	x"07050725",	x"0745072c",	x"07290734",	
					x"073d075f",	x"07650760",	x"07570735",	x"07370745",	
					x"07450751",	x"073c074e",	x"074f0753",	x"075b0732",	
					x"073b0740",	x"073d074f",	x"07630734",	x"07520753",	
					x"0740074e",	x"07410757",	x"075d0764",	x"0759075e",	
					x"0759076d",	x"074f076e",	x"075a0702",	x"112b202f",	
					x"070f0738",	x"071c072c",	x"0745071f",	x"0733071d",	
					x"071906fd",	x"06f00704",	x"070e06d4",	x"06de06b2",	
					x"06de06dd",	x"070b071d",	x"070e0711",	x"070a06fd",	
					x"07080726",	x"073e071f",	x"070c0724",	x"072a06f7",	
					x"07090737",	x"07480757",	x"0730072f",	x"0742071f",	
					x"0715074c",	x"07420755",	x"07390741",	x"073d070b",	
					x"072d0738",	x"072f072d",	x"07300723",	x"0737073b",	
					x"071e0756",	x"07310750",	x"07470755",	x"075006f3",	
					x"112b302f",	x"06f90728",	x"06ef0715",	x"06ec072a",	
					x"0719070c",	x"06ed0706",	x"06f506f6",	x"06f1070b",	
					x"06df06de",	x"06b806e2",	x"070e06e1",	x"06cc0712",	
					x"07100721",	x"0707071b",	x"07400757",	x"0762071a",	
					x"070d0720",	x"06fa0729",	x"07260727",	x"071b072d",	
					x"07410754",	x"0743074e",	x"07400752",	x"073d0750",	
					x"0724071b",	x"070f074d",	x"07260744",	x"0715073d",	
					x"072f0762",	x"07320768",	x"073a0772",	x"07300773",	
					x"074f070c",	x"000a0004",	x"61563ae7",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"112c402f",	x"06ee0714",	x"07150739",	
					x"070e0730",	x"0711070d",	x"06fe073d",	x"06fb072a",	
					x"06fc0705",	x"06ca06e7",	x"06d30714",	x"06e4071b",	
					x"071b072e",	x"0712076b",	x"07240763",	x"0765075e",	
					x"074d0760",	x"075b0747",	x"074a0779",	x"075c0777",	
					x"07700789",	x"076b0775",	x"076b078c",	x"075407a1",	
					x"07730772",	x"07510769",	x"07580787",	x"07640783",	
					x"076b0785",	x"077907bb",	x"075b079e",	x"077307b2",	
					x"078707a1",	x"07820746",	x"112c502f",	x"07210757",	
					x"074e0758",	x"074c0757",	x"07570756",	x"07230744",	
					x"073e074a",	x"07300751",	x"07190723",	x"070a0759",	
					x"073f0774",	x"07520779",	x"07600792",	x"077007a1",	
					x"077d0792",	x"07820799",	x"0772079f",	x"07410792",	
					x"077207a4",	x"078d07ab",	x"079c07c4",	x"07b907d1",	
					x"076907ce",	x"077907b5",	x"0786079a",	x"077607bf",	
					x"078107cf",	x"077d07cc",	x"077e07db",	x"079007d4",	
					x"078607c8",	x"078b07cf",	x"07aa074e",	x"112c602f",	
					x"07040762",	x"07280768",	x"07270778",	x"071e0771",	
					x"072d077e",	x"07580787",	x"07170747",	x"0719072c",	
					x"06e30767",	x"06f207a4",	x"070607b0",	x"078b07dd",	
					x"077b07cc",	x"078807ce",	x"07a207b1",	x"07a707bb",	
					x"078807c5",	x"07cb080b",	x"079807d9",	x"078b07fe",	
					x"07cd07f0",	x"07c50801",	x"07ca07e1",	x"079b07e6",	
					x"07b207fc",	x"07b60811",	x"07c807fb",	x"07bc0806",	
					x"07bf0829",	x"07ba0819",	x"07c2080b",	x"07a9077e",	
					x"112c702f",	x"073807a1",	x"077407c1",	x"077207b4",	
					x"07aa07cf",	x"076107d9",	x"07560763",	x"07680788",	
					x"075f0770",	x"074407ca",	x"076407b6",	x"076e07d6",	
					x"07a30802",	x"07cc080b",	x"07df0816",	x"07d1081c",	
					x"07f90804",	x"07be0837",	x"07f00830",	x"07de0845",	
					x"07f40851",	x"08110835",	x"08070847",	x"08170860",	
					x"081907fd",	x"080d0864",	x"08420874",	x"083e084f",	
					x"0845084d",	x"0820088e",	x"084b086b",	x"083c0870",	
					x"084f06f5",	x"000a0004",	x"85fc7599",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"212d002f",	x"07050707",	x"070706ec",	
					x"06f506ee",	x"06db06f9",	x"06e706da",	x"06bc06b9",	
					x"06d006c9",	x"06bc068f",	x"06a606b0",	x"06ba06cb",	
					x"06d806cc",	x"07030700",	x"06f206f9",	x"06e0071c",	
					x"070c06f3",	x"06f706c4",	x"06eb06f7",	x"071106f9",	
					x"06ee0709",	x"06f006ff",	x"06e60705",	x"070206fd",	
					x"06fc0704",	x"06fe06b6",	x"06c40706",	x"0709071b",	
					x"07190725",	x"06fd0711",	x"07130708",	x"07070731",	
					x"07200730",	x"071506aa",	x"212d102f",	x"06ba06c7",	
					x"06e106ca",	x"06de06fc",	x"06e106fc",	x"06cb06d2",	
					x"06ab06a9",	x"068a0687",	x"067f065f",	x"066b06bb",	
					x"06ad06da",	x"06b106e5",	x"06d206f5",	x"06fa06f9",	
					x"06fe0703",	x"071206d1",	x"06f806cd",	x"06c106d8",	
					x"06e306eb",	x"06e606fb",	x"070506f7",	x"071006f3",	
					x"07080711",	x"07080716",	x"06f306c9",	x"06eb06f0",	
					x"06fe06f2",	x"06e30701",	x"070206ef",	x"06f60704",	
					x"070e0714",	x"07010709",	x"06ec06be",	x"212d202f",	
					x"06c506be",	x"06cb0694",	x"06a106dd",	x"06e106e1",	
					x"06d006b4",	x"06aa0684",	x"066d0680",	x"067d0635",	
					x"066f06b2",	x"06cf06b2",	x"06cc06cd",	x"06e506cc",	
					x"06c306de",	x"06db0701",	x"06db06d6",	x"06d806be",	
					x"06c506cc",	x"06ce06d8",	x"06c306d6",	x"06d406e1",	
					x"06db06c6",	x"06dc06f7",	x"06de06d5",	x"06c906d3",	
					x"06d806e2",	x"06d906df",	x"06c806d5",	x"06eb06e4",	
					x"06c806f7",	x"06ea0713",	x"06f30702",	x"06ef06a6",	
					x"212d302f",	x"069c06a4",	x"069e06c5",	x"069e06af",	
					x"069806d7",	x"069606bd",	x"06890690",	x"06920689",	
					x"066e068c",	x"066b06aa",	x"069406ba",	x"06bd06cb",	
					x"06aa06d0",	x"06ab06d2",	x"06d106ed",	x"06c906d7",	
					x"06bb06ab",	x"069c06da",	x"06c906e9",	x"06cf06f3",	
					x"06cf06e6",	x"06d306ee",	x"070606fa",	x"06e40702",	
					x"06d806bc",	x"06da0718",	x"06ed06de",	x"06d406e4",	
					x"06cb06ee",	x"06ce0724",	x"06fc0722",	x"06fd0726",	
					x"06f6069f",	x"000a0004",	x"73690dc9",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"212e402f",	x"069706ce",	x"06b606e5",	
					x"06c606e0",	x"06d906e3",	x"06cc06ca",	x"06a60699",	
					x"069e06a3",	x"06910685",	x"069506c6",	x"06c806e7",	
					x"06dc0713",	x"071f0723",	x"06e70706",	x"070006fb",	
					x"070a06ff",	x"070f06f5",	x"06fa0709",	x"071f071d",	
					x"070b0733",	x"071c0721",	x"07280737",	x"0715072d",	
					x"0719073e",	x"070e070d",	x"07080742",	x"073d072f",	
					x"070e073f",	x"0727075d",	x"0726076c",	x"07470774",	
					x"072f076b",	x"071c06dc",	x"212e502f",	x"06db0713",	
					x"06fc070d",	x"06e50718",	x"0722071a",	x"06c506eb",	
					x"06d206e7",	x"06bc06ee",	x"06bd06c3",	x"06af071f",	
					x"07140741",	x"07070715",	x"072b0753",	x"0725074e",	
					x"074a0757",	x"07270761",	x"072e071e",	x"070e0752",	
					x"074b074d",	x"071d0751",	x"0744076e",	x"074a076c",	
					x"073f0776",	x"07360762",	x"0735073b",	x"0731076c",	
					x"07430751",	x"071d076a",	x"0734077d",	x"073d0792",	
					x"07470794",	x"07410799",	x"0747070b",	x"212e602f",	
					x"06cc06fe",	x"06ea070d",	x"06ac06fe",	x"06e70701",	
					x"06ea0716",	x"06c8072a",	x"06a00716",	x"06d00713",	
					x"06cd0755",	x"070a074a",	x"07150743",	x"072f078a",	
					x"07440794",	x"07530776",	x"072f0768",	x"0741076c",	
					x"07440783",	x"076a078f",	x"072f077c",	x"075a07a1",	
					x"07670799",	x"076607a0",	x"07550784",	x"0742078c",	
					x"075e079f",	x"074b078a",	x"075707ad",	x"076d07b4",	
					x"076a07cf",	x"077307d0",	x"077d07ca",	x"0792070f",	
					x"212e702f",	x"06e8072a",	x"070e073f",	x"0715075f",	
					x"07210748",	x"070e0725",	x"0730073c",	x"06d4073b",	
					x"06e0071a",	x"06ee07aa",	x"06fb0786",	x"07390791",	
					x"077207a7",	x"077b07a5",	x"077407c2",	x"07b507c1",	
					x"076e07ad",	x"07a207f1",	x"078f07de",	x"078e07ee",	
					x"07a007ed",	x"07c50806",	x"07d307ed",	x"07b6080e",	
					x"07b707cf",	x"079e07f1",	x"07ca07e1",	x"07a307f0",	
					x"07d107f9",	x"07cb082c",	x"07d70843",	x"08090813",	
					x"07e20711",	x"000a0004",	x"9e9b4bdc",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"312f002f",	x"072f073a",	x"0748073f",	
					x"07380752",	x"074a074a",	x"072e0723",	x"07120735",	
					x"071d0730",	x"06e506dd",	x"06d206f6",	x"070f0717",	
					x"071f071b",	x"072c0737",	x"075b0723",	x"0757073e",	
					x"07470758",	x"075d0725",	x"072a073e",	x"07690764",	
					x"074b0733",	x"07520760",	x"0739072d",	x"0739073b",	
					x"0755073a",	x"07290734",	x"07590756",	x"075c073c",	
					x"072d0744",	x"07460746",	x"07330756",	x"07520754",	
					x"07290743",	x"073d0711",	x"312f102f",	x"06f70709",	
					x"0742073a",	x"07350711",	x"072d071d",	x"06f806f4",	
					x"06f60701",	x"06ef06ee",	x"06f006ad",	x"069c0701",	
					x"06e90705",	x"070d0702",	x"07130712",	x"072f072d",	
					x"0751073e",	x"07500727",	x"073806dd",	x"07400716",	
					x"07510739",	x"072f0722",	x"072c074c",	x"073b072e",	
					x"073d0732",	x"07390746",	x"0736071e",	x"074a073e",	
					x"072d0734",	x"072b0726",	x"07320736",	x"071b072a",	
					x"073a073e",	x"0752076b",	x"074d06d2",	x"312f202f",	
					x"06e606f0",	x"071f06f7",	x"07140713",	x"071106f8",	
					x"06ef06f4",	x"06f706d6",	x"06ed06d1",	x"06f606b0",	
					x"069706c4",	x"06e606ee",	x"07210704",	x"06fb06fe",	
					x"06fa0709",	x"072c06ea",	x"06fd073e",	x"072806ed",	
					x"07040714",	x"07140718",	x"072c06fa",	x"06fd071e",	
					x"071e0728",	x"07200727",	x"07140719",	x"071f072e",	
					x"071d074e",	x"072d072b",	x"07370720",	x"0714072c",	
					x"07220725",	x"071c0757",	x"07160748",	x"071206c6",	
					x"312f302f",	x"06cb06e3",	x"06d606f1",	x"06d906f8",	
					x"06e406ea",	x"06cf06f6",	x"06ce06f4",	x"06b706a7",	
					x"06b80695",	x"068b06e8",	x"06df06e8",	x"06d806fc",	
					x"06d80702",	x"06e50712",	x"07150703",	x"06f60701",	
					x"070006d5",	x"06e0070d",	x"07100715",	x"07110724",	
					x"071e071d",	x"072a073c",	x"07350739",	x"071b0711",	
					x"06fe072c",	x"0724073c",	x"072b0721",	x"06ee072f",	
					x"07160720",	x"07000741",	x"071d0757",	x"0726074e",	
					x"071e06e2",	x"000a0004",	x"d48e2c48",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3130402f",	x"06e80703",	x"0700070a",	
					x"06bb070d",	x"07080719",	x"06de06f6",	x"06ea06f8",	
					x"06ec06f8",	x"070206d0",	x"06a906fd",	x"06da072f",	
					x"06e40721",	x"07180737",	x"070e0746",	x"073c0740",	
					x"07380743",	x"07270749",	x"0702075d",	x"0752077e",	
					x"075b0753",	x"0754076a",	x"0741076a",	x"074d075a",	
					x"07580772",	x"0752075d",	x"07460769",	x"07450756",	
					x"074f076d",	x"07630770",	x"074a0798",	x"076b0794",	
					x"07730792",	x"07640713",	x"3130502f",	x"06ef071f",	
					x"07380750",	x"0738074b",	x"073f0737",	x"07150757",	
					x"07150735",	x"071d0720",	x"06f5070b",	x"06fc0767",	
					x"07170768",	x"072a0789",	x"075e0783",	x"073f0789",	
					x"074b07ad",	x"07450792",	x"0732075e",	x"074a07a5",	
					x"077f0795",	x"0747078c",	x"0789079b",	x"0765078f",	
					x"07690793",	x"0761079d",	x"0750079c",	x"077c07bc",	
					x"076e07be",	x"075707c3",	x"078007cd",	x"077207a8",	
					x"078f07f3",	x"079007c0",	x"078f0727",	x"3130602f",	
					x"06fa075e",	x"070f0756",	x"07250772",	x"07550750",	
					x"071f0744",	x"072c0740",	x"070b0731",	x"06eb0736",	
					x"0700076f",	x"06fc077e",	x"0744079c",	x"074807ba",	
					x"078607ae",	x"0780078b",	x"076e07a5",	x"077a077d",	
					x"076b07b9",	x"078f07a5",	x"079207b1",	x"07a607f9",	
					x"078007ba",	x"079707e4",	x"079f07ce",	x"07af07bd",	
					x"079307d1",	x"07ba07e0",	x"078e07dd",	x"07aa07fd",	
					x"079607fd",	x"07a107ed",	x"07a6082b",	x"079f0743",	
					x"3130702f",	x"07230799",	x"076f079e",	x"07870780",	
					x"076d07c2",	x"073c0774",	x"074e0771",	x"074a077f",	
					x"07550771",	x"073f07c5",	x"074a07a7",	x"076507ef",	
					x"079a0826",	x"07ba07f6",	x"07a807ee",	x"07a307fb",	
					x"07d40801",	x"07da080c",	x"07db080d",	x"07d60829",	
					x"07f5084e",	x"07e10828",	x"07ff084c",	x"0811082e",	
					x"081a082c",	x"07f0083b",	x"07fa0850",	x"07fd0842",	
					x"08110859",	x"08150862",	x"08330874",	x"083a088c",	
					x"0823065d",	x"000a0004",	x"fab669a5",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"01310030",	x"068f066a",	x"0656065a",	
					x"0663065a",	x"06620645",	x"06380659",	x"0642068b",	
					x"0695069f",	x"06d20655",	x"0664068c",	x"06bd06bb",	
					x"06b006b0",	x"06960690",	x"06940692",	x"068c0682",	
					x"068a0694",	x"068d062a",	x"065b0666",	x"06960699",	
					x"0691068a",	x"06930695",	x"069b06a0",	x"068e069a",	
					x"06b5069e",	x"06980661",	x"06670687",	x"06af06a9",	
					x"06ab06a5",	x"06b2069f",	x"069c06a7",	x"069706d1",	
					x"06a00691",	x"0681064a",	x"01311030",	x"065a0637",	
					x"063a0631",	x"06310634",	x"065e061c",	x"06210656",	
					x"063e067b",	x"06600679",	x"0672064b",	x"066f0647",	
					x"067d0685",	x"068c0685",	x"06860655",	x"068d0680",	
					x"069f0695",	x"06a3068f",	x"069e0615",	x"06680673",	
					x"068e066e",	x"0672065b",	x"06890681",	x"0679068f",	
					x"068a067c",	x"06750674",	x"06910644",	x"06870678",	
					x"0691067c",	x"0690068b",	x"0687068c",	x"068f0690",	
					x"06b00697",	x"0697067e",	x"06790637",	x"01312030",	
					x"064c0647",	x"063c0657",	x"06450607",	x"061e0618",	
					x"06440629",	x"06730665",	x"067f064f",	x"066d063a",	
					x"064f063e",	x"0656063d",	x"0660064d",	x"0651065e",	
					x"067e0664",	x"06740669",	x"066a0659",	x"0675063f",	
					x"0665065d",	x"065e064e",	x"064c0643",	x"066e0647",	
					x"0663064d",	x"064b0681",	x"06870677",	x"06560639",	
					x"06530670",	x"066b0672",	x"067a0673",	x"067d0681",	
					x"066c064b",	x"06650685",	x"0663065d",	x"065e062d",	
					x"01313030",	x"0634063e",	x"0615061b",	x"0607061c",	
					x"06210618",	x"06090632",	x"06380654",	x"0650064f",	
					x"0645061e",	x"063b0636",	x"0644065c",	x"064d065c",	
					x"06660659",	x"06590657",	x"0662067c",	x"066d0660",	
					x"06550628",	x"0632063d",	x"064b0649",	x"0653063e",	
					x"0655065e",	x"065b0674",	x"06760691",	x"0682066b",	
					x"065b0622",	x"0642066e",	x"066f067f",	x"0660067a",	
					x"06700691",	x"066b0699",	x"06760695",	x"06650680",	
					x"06820628",	x"000a0004",	x"bf7ad247",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"01324030",	x"064d063a",	x"06320629",	
					x"06000620",	x"06220634",	x"060d062f",	x"064f0659",	
					x"0665066f",	x"0640064d",	x"063d0671",	x"065e066b",	
					x"065b0681",	x"069b0678",	x"0662067b",	x"067c0689",	
					x"0691068d",	x"06890649",	x"0650069c",	x"0668067e",	
					x"06970686",	x"067f0693",	x"06a006a0",	x"069b069c",	
					x"069e0687",	x"06960676",	x"06860697",	x"069806b7",	
					x"06a106b7",	x"06bd06bc",	x"069d06be",	x"06b406ba",	
					x"06a706b3",	x"06ba067a",	x"01325030",	x"066e0670",	
					x"065d0667",	x"064c0663",	x"0678068a",	x"0684068a",	
					x"06830685",	x"068a068f",	x"06960687",	x"06840698",	
					x"069206be",	x"069106a8",	x"06a206be",	x"06b806b8",	
					x"06b706b7",	x"06b506b7",	x"069f06b2",	x"068c06a7",	
					x"06aa06a9",	x"069e06b1",	x"06b806c0",	x"06b906d4",	
					x"06b006c0",	x"06b106b2",	x"069e06a6",	x"06a506e8",	
					x"06bb06c9",	x"06cb06f0",	x"06cd0704",	x"06c506e8",	
					x"06ba06e9",	x"06cf06cd",	x"06c00693",	x"01326030",	
					x"069706a0",	x"06740690",	x"067b0692",	x"068406a0",	
					x"067506af",	x"06940697",	x"0694069f",	x"06a1069f",	
					x"067c0699",	x"068106ec",	x"06c206be",	x"06c906e6",	
					x"06e606f8",	x"06e006db",	x"06e706d0",	x"06cb06cc",	
					x"06b206e1",	x"06cf06d8",	x"06d406ef",	x"06ec0709",	
					x"06e90703",	x"06ea070c",	x"06fe06fc",	x"06c906d0",	
					x"06d00714",	x"0704070c",	x"0700070c",	x"06fe0718",	
					x"06f60716",	x"06f0073a",	x"06f8072f",	x"070a06d5",	
					x"01327030",	x"06c1070b",	x"068506c6",	x"068e069f",	
					x"06a506d9",	x"06bb06e2",	x"06e20708",	x"06f906ee",	
					x"06bd06d7",	x"06d30723",	x"0719072b",	x"07210718",	
					x"07150746",	x"072c0765",	x"0748075b",	x"073b0739",	
					x"073a0704",	x"07080743",	x"073e0733",	x"0722074a",	
					x"07420778",	x"076f0787",	x"077b077b",	x"076e0746",	
					x"075f0744",	x"0760076f",	x"0770079c",	x"07710780",	
					x"079307b5",	x"077a07a1",	x"077b07b4",	x"07880781",	
					x"07790720",	x"000a0004",	x"e9390855",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"11330030",	x"07450709",	x"06ee0716",	
					x"07220705",	x"072a0707",	x"06ff070e",	x"0713071a",	
					x"071f0720",	x"073d070f",	x"072f0764",	x"076b075f",	
					x"07700760",	x"0771074e",	x"0773072e",	x"0753073f",	
					x"074b0739",	x"07760710",	x"07470733",	x"0761074c",	
					x"0751073b",	x"075d0760",	x"07500746",	x"0735075d",	
					x"0754073a",	x"073406fa",	x"06fc075d",	x"07520747",	
					x"07480752",	x"074c0769",	x"0744073c",	x"07610777",	
					x"074f0749",	x"073c0718",	x"11331030",	x"06f706ff",	
					x"07200704",	x"070906e4",	x"070b06fc",	x"06e70702",	
					x"06f70703",	x"07100720",	x"072b0707",	x"073a073c",	
					x"07370737",	x"072e0736",	x"07470735",	x"072e0737",	
					x"07340739",	x"07530758",	x"076f070d",	x"07380720",	
					x"074c0743",	x"0745074d",	x"075e071b",	x"07400732",	
					x"072d0732",	x"07250741",	x"0736071e",	x"0740074d",	
					x"073f075a",	x"074e0761",	x"07530755",	x"073e074f",	
					x"0754074a",	x"0730076a",	x"074606e1",	x"11332030",	
					x"070606dd",	x"06f606e2",	x"070606f0",	x"070d06fc",	
					x"071406fe",	x"0711071b",	x"07300730",	x"073d0713",	
					x"072c0719",	x"07530731",	x"072f0730",	x"071a0705",	
					x"07150712",	x"07240728",	x"0732072c",	x"07450703",	
					x"06fe071c",	x"07260728",	x"0719071e",	x"07150716",	
					x"07110725",	x"0736073c",	x"071c071e",	x"07180705",	
					x"07170729",	x"0755072a",	x"07310741",	x"074c0751",	
					x"0737074f",	x"073c0742",	x"0716073d",	x"073306e8",	
					x"11333030",	x"06d806cf",	x"06d606df",	x"06d806dd",	
					x"06dc06f6",	x"06e406e4",	x"06e706d6",	x"06e406fc",	
					x"06e106cc",	x"06ea0709",	x"0705072a",	x"0719072a",	
					x"071f06f2",	x"06f90712",	x"07130733",	x"072b0714",	
					x"07190713",	x"07160738",	x"07220726",	x"071f0717",	
					x"07220712",	x"070d0712",	x"07080718",	x"071a0740",	
					x"072f071c",	x"071b074e",	x"075b074a",	x"073c0745",	
					x"07350745",	x"0724074b",	x"0728074d",	x"07220744",	
					x"072706ee",	x"000a0004",	x"5dcb3277",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"11344030",	x"06fb06f0",	x"06e606f8",	
					x"06d2070a",	x"070a0709",	x"07000725",	x"071c072b",	
					x"07230723",	x"07350702",	x"0704071e",	x"07180744",	
					x"0733074b",	x"07390755",	x"07410742",	x"073f0744",	
					x"07520743",	x"07370732",	x"0740077b",	x"0749074c",	
					x"0741076b",	x"075f0749",	x"07440759",	x"07520759",	
					x"0756076f",	x"0762075e",	x"075b0774",	x"07680774",	
					x"077e0779",	x"077e0788",	x"0779078d",	x"077b079d",	
					x"07700783",	x"076a0730",	x"11345030",	x"0738072b",	
					x"07330728",	x"0723073e",	x"07250752",	x"074c0739",	
					x"075f0776",	x"07530751",	x"074d0748",	x"07480783",	
					x"0778076f",	x"07560765",	x"07740782",	x"07810785",	
					x"0773077a",	x"076b0762",	x"07540766",	x"0756078c",	
					x"0783078b",	x"0780078a",	x"0779078f",	x"076e07b8",	
					x"077907b0",	x"078107a4",	x"0777079e",	x"075f079a",	
					x"078007b1",	x"078107af",	x"077707b7",	x"078907a3",	
					x"077c07c5",	x"078e07c4",	x"0797072c",	x"11346030",	
					x"06f40749",	x"0728074d",	x"073d075e",	x"07430760",	
					x"07480748",	x"07360769",	x"077e075f",	x"07510765",	
					x"075b0794",	x"078907a3",	x"078d079e",	x"07a607a7",	
					x"07a807b0",	x"079a07b1",	x"077507b1",	x"079c07ac",	
					x"07a107a7",	x"07c707ba",	x"07ab07ae",	x"07bd07b0",	
					x"07a007b1",	x"07a907c5",	x"07ae07c3",	x"07b007bb",	
					x"078707e3",	x"07c307f8",	x"07cd07ff",	x"07c80800",	
					x"07bf080f",	x"07cf07ea",	x"07ca07d8",	x"07ab07ac",	
					x"11347030",	x"078f07c5",	x"079507af",	x"078a07c8",	
					x"077407dc",	x"078507ac",	x"079307d6",	x"07bc07d8",	
					x"07d507ee",	x"078907f4",	x"07ce0820",	x"07f6081f",	
					x"08070805",	x"07f80805",	x"08160829",	x"0807081f",	
					x"0803080a",	x"07f6081c",	x"08210825",	x"080d0840",	
					x"081d084a",	x"08170845",	x"08300853",	x"08320835",	
					x"08380835",	x"0843084b",	x"08480850",	x"08570850",	
					x"084b0862",	x"084d0879",	x"08430843",	x"083b0868",	
					x"084b06da",	x"000a0004",	x"8e8b6f8b",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"21350030",	x"06e406a7",	x"06a1069e",	
					x"069906cc",	x"06c006bf",	x"06c306ba",	x"06e606ba",	
					x"06e006ba",	x"06e806c4",	x"06c406f0",	x"06eb0701",	
					x"06ed06ec",	x"070906ee",	x"06f50700",	x"06d30710",	
					x"071106f0",	x"070206a0",	x"06d506dc",	x"070306cc",	
					x"0700072c",	x"070206e1",	x"06f206fb",	x"071206ff",	
					x"070206eb",	x"06e806ac",	x"06e00706",	x"070e0725",	
					x"06ff0721",	x"07180720",	x"06f806f5",	x"06e006ff",	
					x"06e806e2",	x"06ed0677",	x"21351030",	x"069206b8",	
					x"06b106a8",	x"06a4067f",	x"069a06b1",	x"06ab06c5",	
					x"06ca06dd",	x"06e906d8",	x"06c506b4",	x"06c306f0",	
					x"06fd0706",	x"06f6070d",	x"06f706e6",	x"06f406e1",	
					x"06d806d6",	x"06f806c3",	x"06f306a9",	x"06d206d7",	
					x"06dd06ce",	x"06ee06e3",	x"06fb06e9",	x"06eb06ed",	
					x"06ff06ed",	x"06f106e1",	x"06ec06a8",	x"06d706f0",	
					x"06ef06f0",	x"06f106f6",	x"06f906ef",	x"06ef0728",	
					x"070706f9",	x"06fb0706",	x"06f20686",	x"21352030",	
					x"06930685",	x"069a06a4",	x"069206a2",	x"06ad069b",	
					x"06b50690",	x"06be06b6",	x"06c806ad",	x"06d506a3",	
					x"06c106cd",	x"06d406e2",	x"06e006eb",	x"06e306de",	
					x"06e206d7",	x"06c806db",	x"06cb06e6",	x"06db069e",	
					x"06a906bd",	x"06c806d8",	x"06ae06ca",	x"06d006c5",	
					x"06d006d4",	x"06d306e7",	x"06f006d8",	x"06b106a2",	
					x"06b206e1",	x"06c706f0",	x"06dd06e7",	x"06f00701",	
					x"06c406ec",	x"06d406f6",	x"06de06e3",	x"06d206ac",	
					x"21353030",	x"069f067a",	x"067306a3",	x"06900682",	
					x"068c06b5",	x"069a06ba",	x"06c006ab",	x"06ae06a8",	
					x"06a60685",	x"069906bd",	x"06b906d9",	x"06da06d5",	
					x"06db06dc",	x"06c106ae",	x"06cb06c8",	x"06bb06db",	
					x"06c3069f",	x"069306d9",	x"06dd06ef",	x"06e606d7",	
					x"06db06d2",	x"06c006d7",	x"06d006da",	x"06cf06e8",	
					x"06c306ab",	x"06bc06ee",	x"06ef0700",	x"06de06e6",	
					x"06d106fd",	x"06d306fa",	x"06d7070a",	x"06d90701",	
					x"06eb0698",	x"000a0004",	x"72f30945",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"21364030",	x"06ac06b0",	x"069006c1",	
					x"06ac06c0",	x"06b506c9",	x"06ba06cf",	x"06c806bc",	
					x"06b506c0",	x"06b606ba",	x"06cd06df",	x"06db06ec",	
					x"070106f1",	x"070c0700",	x"06dc06eb",	x"06d806f5",	
					x"06f106eb",	x"06fc06d7",	x"06d306ff",	x"07140708",	
					x"06ff0700",	x"070f06e9",	x"07090706",	x"0708070b",	
					x"071a0716",	x"07080705",	x"06ed0739",	x"07280708",	
					x"0703072b",	x"07180721",	x"070f0721",	x"07170728",	
					x"071f072b",	x"071a06b9",	x"21365030",	x"06bc06d8",	
					x"06da06e8",	x"06c606df",	x"06d006ee",	x"06d906f2",	
					x"06dd0718",	x"070c0701",	x"07020708",	x"06fe0729",	
					x"0705072c",	x"071f0729",	x"0726073e",	x"070a0717",	
					x"0729072a",	x"07140726",	x"070d0715",	x"070a072a",	
					x"07280730",	x"072e072c",	x"07120755",	x"072f074d",	
					x"0728074c",	x"0719074f",	x"07270733",	x"0722075b",	
					x"07330765",	x"0741077b",	x"07410776",	x"074d077f",	
					x"074a0753",	x"07310757",	x"073a06e9",	x"21366030",	
					x"06d306f8",	x"06f906eb",	x"06cf06f2",	x"06f70718",	
					x"0715071c",	x"071c0723",	x"0717071a",	x"06f0071b",	
					x"07030734",	x"071c073e",	x"07370745",	x"07550762",	
					x"0760075c",	x"07420755",	x"07370750",	x"073e0734",	
					x"07230757",	x"07550798",	x"07570761",	x"075d075d",	
					x"075b0756",	x"07350780",	x"074b0761",	x"074e075f",	
					x"074d0787",	x"076007b2",	x"0762078c",	x"0773079f",	
					x"0774079c",	x"077007a7",	x"0775079e",	x"07750722",	
					x"21367030",	x"072c0772",	x"071c0727",	x"07100747",	
					x"073a0773",	x"074d076d",	x"07540769",	x"076b0776",	
					x"07380773",	x"07430792",	x"077507c4",	x"079907ad",	
					x"07a707bb",	x"07a807b6",	x"07a107f3",	x"07a807c7",	
					x"079907ac",	x"07ba07d4",	x"07e607da",	x"07c707d3",	
					x"07d507d0",	x"07d707e1",	x"07d307c5",	x"07ca07dd",	
					x"07d007de",	x"07d907f9",	x"07e807e4",	x"07ea080a",	
					x"07ee0816",	x"07f1080f",	x"07f40824",	x"07f5080e",	
					x"07fd06dd",	x"000a0004",	x"a4464472",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"31370030",	x"06fb0705",	x"071006fc",	
					x"06f206d9",	x"06fa06fc",	x"071d072b",	x"070a0723",	
					x"07100718",	x"07170705",	x"073e0738",	x"076c0753",	
					x"0751071b",	x"07430743",	x"0757073f",	x"074a0721",	
					x"07320723",	x"071a06d3",	x"07180726",	x"07390738",	
					x"0744072d",	x"0745072c",	x"07340747",	x"07390731",	
					x"072d071c",	x"072b06f7",	x"06fd0723",	x"07530755",	
					x"0753075e",	x"077a0750",	x"075c0734",	x"07440742",	
					x"071b0719",	x"071a06b0",	x"31371030",	x"06e006a9",	
					x"06d806fc",	x"06e406c2",	x"06db06cb",	x"06ea0700",	
					x"07170706",	x"0715070c",	x"071206ce",	x"06f80719",	
					x"0724073e",	x"073b071d",	x"0756075a",	x"073d0708",	
					x"07290733",	x"0711072c",	x"071606da",	x"06f1070f",	
					x"07220715",	x"07220738",	x"074f073c",	x"072b072f",	
					x"07210712",	x"071206f9",	x"070806fd",	x"06fd071c",	
					x"07110725",	x"07350738",	x"07450748",	x"07420737",	
					x"073c071f",	x"0725073c",	x"072206da",	x"31372030",	
					x"071806b3",	x"06d206c1",	x"06ff06bc",	x"06e506d2",	
					x"06f3071a",	x"06f806de",	x"070306f2",	x"070f06bc",	
					x"06fb0704",	x"07340711",	x"072c072d",	x"072c06f8",	
					x"071406fb",	x"071806f6",	x"06f306fb",	x"06fe06d0",	
					x"06f90708",	x"071c0710",	x"072b0721",	x"07100711",	
					x"0718072b",	x"0716071b",	x"0708070d",	x"06fa06dd",	
					x"06ee071d",	x"070c0716",	x"0726071f",	x"071e071b",	
					x"0706071b",	x"07170724",	x"06fb072c",	x"06f806bb",	
					x"31373030",	x"06c806c0",	x"06cf06a1",	x"06ba06b4",	
					x"06c906ac",	x"06ae06c9",	x"06d906ed",	x"06cc06dd",	
					x"06e606c1",	x"06d606e8",	x"06ef06fd",	x"07040719",	
					x"07060706",	x"06e20707",	x"06ff0717",	x"070306f4",	
					x"06ea0697",	x"06c206f7",	x"06fe070e",	x"06f9071c",	
					x"07200711",	x"070a06fb",	x"06f4070c",	x"06f30705",	
					x"06ff06f5",	x"06fc071c",	x"07170717",	x"070d071a",	
					x"071b072f",	x"0722071c",	x"07150716",	x"0705071d",	
					x"070b06c9",	x"000a0004",	x"d1542414",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"31384030",	x"06f706d4",	x"06c706d8",	
					x"06cb06d6",	x"06da06e2",	x"06d206ed",	x"06dd071d",	
					x"070f06f5",	x"070406ff",	x"070f0716",	x"072d0746",	
					x"0725071e",	x"07380726",	x"070e072f",	x"073d0728",	
					x"07090711",	x"071c0709",	x"06f90730",	x"073e072c",	
					x"072c074c",	x"07530756",	x"073a0724",	x"07340742",	
					x"07390745",	x"073b072d",	x"072f0741",	x"07420763",	
					x"07620773",	x"07730777",	x"07630766",	x"0762076b",	
					x"0761075a",	x"0752070f",	x"31385030",	x"070a0721",	
					x"06f5072a",	x"0715072b",	x"07310732",	x"0718074c",	
					x"07310746",	x"073e0735",	x"072e073c",	x"07400764",	
					x"07520763",	x"07530763",	x"07630777",	x"07590763",	
					x"075e077b",	x"074c075e",	x"074a0741",	x"07280771",	
					x"0773077c",	x"07540776",	x"07710789",	x"075f076e",	
					x"07620775",	x"0737078d",	x"0747076c",	x"073b07a7",	
					x"076a07af",	x"077907a7",	x"077e07ae",	x"077f079b",	
					x"076707a3",	x"076f0792",	x"07490726",	x"31386030",	
					x"06f80746",	x"07030750",	x"07280704",	x"070c075b",	
					x"073e0766",	x"073e075d",	x"07590750",	x"07420738",	
					x"0735076c",	x"0749079d",	x"076a079f",	x"07770793",	
					x"078f078e",	x"076a0787",	x"07570788",	x"07600768",	
					x"077207a8",	x"07a107b5",	x"079107a6",	x"07ad07c7",	
					x"079607a2",	x"079407ab",	x"079207a8",	x"079d07ab",	
					x"079307d7",	x"07b707e0",	x"07a407cf",	x"07ac07e5",	
					x"079307cb",	x"078a07c3",	x"079407db",	x"079e0775",	
					x"31387030",	x"076a0795",	x"0782079d",	x"07960797",	
					x"07710785",	x"07520767",	x"076307b1",	x"07b407b2",	
					x"07be07a2",	x"07920803",	x"07df0800",	x"07f50810",	
					x"07e90816",	x"07eb080a",	x"07f607f4",	x"07d60806",	
					x"07ec07df",	x"07e80802",	x"080e0814",	x"0800081e",	
					x"080d0840",	x"0829081f",	x"081b081d",	x"07e60818",	
					x"082c0832",	x"08270839",	x"082d0841",	x"08260845",	
					x"08440878",	x"08200881",	x"08380872",	x"083d0846",	
					x"08280660",	x"000a0004",	x"018462a2",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"01390031",	x"0690065f",	x"06580664",	
					x"0668064a",	x"06440648",	x"06420653",	x"063a0643",	
					x"063e0645",	x"06470634",	x"062b066d",	x"064e0696",	
					x"067a0699",	x"06b60691",	x"06710668",	x"067d0675",	
					x"065f0669",	x"06760645",	x"06510666",	x"06750692",	
					x"0688066b",	x"06970689",	x"06740695",	x"0688068a",	
					x"068d0667",	x"06850655",	x"06630686",	x"06880678",	
					x"067f0679",	x"06750689",	x"06820687",	x"068706cb",	
					x"068e067e",	x"0670062d",	x"01391031",	x"066f0633",	
					x"0653065a",	x"06590633",	x"06450639",	x"063b0628",	
					x"06210630",	x"0619061b",	x"0628062d",	x"064a0660",	
					x"0658067b",	x"066a067f",	x"06820664",	x"067f0669",	
					x"067d0667",	x"06700667",	x"066e0630",	x"063d068b",	
					x"06800652",	x"066c0671",	x"06890685",	x"068c067d",	
					x"067c0672",	x"0663066b",	x"06710658",	x"06670656",	
					x"06940694",	x"06a10694",	x"0697068d",	x"06860689",	
					x"06980694",	x"068d0688",	x"0687063c",	x"01392031",	
					x"06320635",	x"06410665",	x"064c0629",	x"06230626",	
					x"0638061a",	x"064a0646",	x"06500649",	x"06590617",	
					x"064b0636",	x"06620662",	x"06730681",	x"0672066c",	
					x"0673064f",	x"06720649",	x"064c0654",	x"06590632",	
					x"06630654",	x"06630663",	x"065d065d",	x"06810661",	
					x"0662066c",	x"065e0668",	x"065b0661",	x"065b0653",	
					x"065c0672",	x"0660067c",	x"066d0679",	x"06940678",	
					x"0681065e",	x"067d0675",	x"066f067d",	x"06750622",	
					x"01393031",	x"063e0642",	x"061d063c",	x"061b0628",	
					x"061e0625",	x"060c061e",	x"0619061f",	x"061a0632",	
					x"06320621",	x"0627065e",	x"06510662",	x"064f065d",	
					x"0670065c",	x"06450642",	x"0649066b",	x"06570657",	
					x"06540651",	x"064f0654",	x"064e0671",	x"06550669",	
					x"066d0675",	x"064a0683",	x"0670068a",	x"0677067a",	
					x"0651065f",	x"064c066e",	x"064c0683",	x"06690692",	
					x"067e0693",	x"066d06a1",	x"066906a7",	x"066f068d",	
					x"0670062b",	x"000a0004",	x"b970d011",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"013a4031",	x"063d0626",	x"062f0649",	
					x"064a0639",	x"06370631",	x"06030645",	x"06390648",	
					x"063f0668",	x"063f062e",	x"06300667",	x"0643067b",	
					x"06640688",	x"06910679",	x"06710685",	x"067a0683",	
					x"068706a1",	x"0673066a",	x"066c06c1",	x"06ac06b7",	
					x"069c0699",	x"06a506c3",	x"069206c3",	x"06c106bb",	
					x"0691068f",	x"069b069c",	x"068f06bb",	x"06a106cf",	
					x"06b406d6",	x"06cb06d3",	x"06c906e0",	x"06c706de",	
					x"06b706b9",	x"06b1065b",	x"013a5031",	x"066b068a",	
					x"06730692",	x"0683067a",	x"067a067f",	x"06560693",	
					x"066d0690",	x"067906a6",	x"068c06a2",	x"067e06b4",	
					x"06af06c1",	x"06bc06d2",	x"06ce06f5",	x"06a606b6",	
					x"06b006c8",	x"06af06cb",	x"069c06bd",	x"06a406e6",	
					x"06a806dd",	x"06a006e5",	x"06c206dd",	x"06c106fd",	
					x"06c406e7",	x"06c006dc",	x"06ae06ca",	x"06ae06fc",	
					x"06c806f2",	x"06c106e3",	x"06ad070b",	x"06d00704",	
					x"06d30709",	x"06de06e4",	x"06c90691",	x"013a6031",	
					x"067306ae",	x"069006ac",	x"067f069d",	x"067a069e",	
					x"06860693",	x"0687068a",	x"0677068d",	x"065a069e",	
					x"067906e2",	x"06be06e0",	x"06cf06df",	x"06e106e3",	
					x"06d706f7",	x"06d50713",	x"06c80704",	x"06e806ea",	
					x"06e40716",	x"06c406fe",	x"06e80711",	x"06f90717",	
					x"06ee0717",	x"06f5072b",	x"07150742",	x"06f506f2",	
					x"06e00735",	x"06f4072d",	x"06f70749",	x"06ff072e",	
					x"0712074a",	x"07070738",	x"07050730",	x"06f206c5",	
					x"013a7031",	x"06b106f8",	x"06ac0704",	x"06a906c2",	
					x"06a506e3",	x"06a106dd",	x"06bc071f",	x"06dd06f2",	
					x"06d406c8",	x"06c1072f",	x"0720075f",	x"072a073c",	
					x"0720074f",	x"072d074d",	x"071c0761",	x"07340768",	
					x"0734071c",	x"072f0773",	x"07640772",	x"074b0781",	
					x"074a0789",	x"07650794",	x"07600797",	x"077f0787",	
					x"075c076e",	x"075c079d",	x"076507c6",	x"078e07a2",	
					x"07a807cd",	x"07af07a1",	x"077a07cd",	x"0782079e",	
					x"07910717",	x"000a0004",	x"ec121344",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"113b0031",	x"0753074f",	x"0772074f",	
					x"07650767",	x"077d073f",	x"072e071f",	x"07160722",	
					x"07040726",	x"070306e0",	x"06df0716",	x"072306f1",	
					x"0728072b",	x"073b0739",	x"074b073a",	x"07650770",	
					x"07640725",	x"077a071e",	x"071f074f",	x"07840738",	
					x"073c073d",	x"075d073d",	x"074f073e",	x"07500745",	
					x"0746076f",	x"076106e2",	x"070d0739",	x"07380744",	
					x"07410758",	x"07550761",	x"072e073e",	x"073c0758",	
					x"073a0748",	x"0754072d",	x"113b1031",	x"0739073e",	
					x"0759074b",	x"0752073c",	x"074f0718",	x"070b072e",	
					x"070806e9",	x"06da06fe",	x"06f106cb",	x"06d606e5",	
					x"06ee0702",	x"06f80709",	x"07040717",	x"0748074f",	
					x"07410719",	x"074d0744",	x"0759072b",	x"07260754",	
					x"07600767",	x"074d0748",	x"07520737",	x"07570736",	
					x"074c0759",	x"07500756",	x"0756070e",	x"07140731",	
					x"073e0740",	x"07410738",	x"07500749",	x"0747073d",	
					x"076a0772",	x"075d0777",	x"0748071d",	x"113b2031",	
					x"072c0741",	x"0709071f",	x"0716072e",	x"0737071c",	
					x"07220703",	x"070f06fe",	x"070406f6",	x"06f006ca",	
					x"06f406e3",	x"070306f9",	x"06ef06e9",	x"06fc06f2",	
					x"07170729",	x"0739071d",	x"071a071f",	x"071906f9",	
					x"06f80722",	x"0721074f",	x"0736072c",	x"072c0724",	
					x"071c0740",	x"072b074b",	x"072a0727",	x"071906ef",	
					x"07040733",	x"07290723",	x"072f0722",	x"07400741",	
					x"071c0748",	x"0745074b",	x"07460742",	x"073b06f1",	
					x"113b3031",	x"06eb0715",	x"06ee0702",	x"06e70700",	
					x"071206ff",	x"06f406e4",	x"06d206f8",	x"06df06db",	
					x"06c806e3",	x"06d206ed",	x"06e706ed",	x"06c60706",	
					x"07080732",	x"07160735",	x"072b0745",	x"072e0718",	
					x"070e071a",	x"07070747",	x"072b071c",	x"0725076c",	
					x"073d0743",	x"07370737",	x"0730073f",	x"073c0753",	
					x"072a0725",	x"0715075d",	x"07340751",	x"07220746",	
					x"07360750",	x"07340763",	x"072f0762",	x"0723075c",	
					x"072d0717",	x"000a0004",	x"5d4334e1",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"113c4031",	x"06fb0738",	x"07200746",	
					x"07240728",	x"0716072d",	x"06ec0727",	x"0708071f",	
					x"06f4070a",	x"06cc06d7",	x"06e2070c",	x"06d60716",	
					x"0715072a",	x"072a0769",	x"07140755",	x"0747076b",	
					x"074c0751",	x"073c074f",	x"0749076f",	x"07680792",	
					x"077f0798",	x"07510769",	x"07700785",	x"076a0781",	
					x"0771077d",	x"0764076c",	x"075b07a5",	x"077607b1",	
					x"07640782",	x"07780781",	x"0765079f",	x"078307bc",	
					x"078a07a8",	x"077a0748",	x"113c5031",	x"074d0765",	
					x"074a0772",	x"075a075e",	x"0765078f",	x"0737074f",	
					x"0756073a",	x"07440742",	x"0734073a",	x"07090754",	
					x"07500761",	x"075b0782",	x"07660791",	x"0793079d",	
					x"074f0799",	x"078407a0",	x"076c078b",	x"0753079f",	
					x"078507af",	x"076807a5",	x"077507a2",	x"078b07b6",	
					x"078c07d1",	x"078a07cf",	x"078e07b7",	x"076507c3",	
					x"07a907cc",	x"079207cd",	x"078607d0",	x"079507d0",	
					x"078e07fc",	x"079e07c2",	x"07900751",	x"113c6031",	
					x"074d076d",	x"074e077b",	x"07530781",	x"07680771",	
					x"074b077e",	x"0748077c",	x"07520769",	x"0714073b",	
					x"071d078a",	x"075107b3",	x"0756079b",	x"079307d4",	
					x"07a107bb",	x"079207be",	x"079507d4",	x"077e07bf",	
					x"077e07db",	x"07ad07f2",	x"07b107e0",	x"07c507dc",	
					x"07b107f5",	x"07c007fc",	x"07cc07e0",	x"07b407cd",	
					x"07a607f7",	x"07de07f8",	x"07c0080a",	x"07c107fd",	
					x"07bf0833",	x"07bc080c",	x"07ac0819",	x"07c7079a",	
					x"113c7031",	x"078a07bb",	x"079b07bb",	x"079207d0",	
					x"079907d8",	x"07a207bd",	x"07a007ca",	x"07a507a2",	
					x"079c079a",	x"077507e2",	x"078e07cc",	x"07b10813",	
					x"07b20817",	x"07e5082b",	x"08150837",	x"07f50838",	
					x"08010840",	x"07cb086a",	x"082a0863",	x"082f0872",	
					x"08290876",	x"083b0857",	x"08360862",	x"08480889",	
					x"082f0844",	x"08410858",	x"085b086e",	x"0858086a",	
					x"085b085e",	x"0850089c",	x"086c08a2",	x"0877088b",	
					x"085706c7",	x"000a0004",	x"8ed67a0e",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"213d0031",	x"06dd06e2",	x"070706e3",	
					x"06e906f2",	x"06e5070a",	x"06e906a5",	x"06b106b7",	
					x"06c506a8",	x"0698067e",	x"0684069a",	x"06c806b3",	
					x"06e306eb",	x"070d0703",	x"071506fa",	x"07010702",	
					x"070a06ea",	x"06f706ab",	x"06d006e1",	x"06f506e7",	
					x"06f506f8",	x"070606ee",	x"06f906f4",	x"06f306df",	
					x"06e50705",	x"06db06b7",	x"06da06e6",	x"070806ee",	
					x"06e406f3",	x"06ef06f8",	x"06ea0710",	x"06f6072b",	
					x"0716071a",	x"071606be",	x"213d1031",	x"06d206c6",	
					x"06da06d7",	x"06cc06ce",	x"06dd06cb",	x"06c606c1",	
					x"06a806bb",	x"067d0678",	x"06580650",	x"06730675",	
					x"066706bd",	x"06a606be",	x"06b406d6",	x"06d606c7",	
					x"06de070e",	x"070306c5",	x"06dc0694",	x"069f06d7",	
					x"06e506d6",	x"06de06de",	x"06f106d7",	x"06e506e7",	
					x"06f906e7",	x"06e506eb",	x"06e306b6",	x"06df06e7",	
					x"06d906e2",	x"06d906e8",	x"06e606f8",	x"06e1070a",	
					x"06ee0727",	x"072b070a",	x"06fa06ac",	x"213d2031",	
					x"06e006a9",	x"06bc06b0",	x"06c606b7",	x"06d806a3",	
					x"06bb0693",	x"06930697",	x"06810692",	x"0688063b",	
					x"066d0689",	x"06a00681",	x"06a306c4",	x"06d506ce",	
					x"06d206ec",	x"06d206cc",	x"06d706bf",	x"06bf06bc",	
					x"06bd06cc",	x"06d206fd",	x"06d706d1",	x"06d106d3",	
					x"06b206cd",	x"06d106df",	x"06e906ed",	x"06d606b9",	
					x"06c406d8",	x"06ca06bf",	x"06c506dc",	x"06f406e9",	
					x"06cf06e8",	x"06df070e",	x"06ed06fc",	x"06f4069c",	
					x"213d3031",	x"069106a3",	x"069306ad",	x"06ae06a9",	
					x"069b06b7",	x"069006af",	x"06970691",	x"068a066c",	
					x"067e065f",	x"0668069a",	x"068c06bd",	x"06c406bc",	
					x"06bd06e4",	x"06ba06d0",	x"06d006d1",	x"06b306e1",	
					x"06b906b5",	x"06a206d7",	x"06bc06f5",	x"06d406e0",	
					x"06ce06de",	x"06c306ed",	x"06dc06dc",	x"06db06db",	
					x"06c206ca",	x"06c30704",	x"06d506cb",	x"06c206e2",	
					x"06ca06f1",	x"06d606ff",	x"06d90721",	x"0704071c",	
					x"06eb06a1",	x"000a0004",	x"6f73070f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"213e4031",	x"06ad06c3",	x"06be06d7",	
					x"06bb06e1",	x"06c106c9",	x"06bf06b6",	x"06aa06a7",	
					x"068d06a2",	x"06b60694",	x"066506d6",	x"06be06e5",	
					x"06f106ef",	x"06fa0711",	x"06ed0700",	x"0701070f",	
					x"07030704",	x"06fc06e3",	x"06d606fb",	x"0716072c",	
					x"0710074e",	x"0712072b",	x"071c0722",	x"0706072c",	
					x"0725072f",	x"07260713",	x"06fc0726",	x"070e0733",	
					x"070d073c",	x"071e0748",	x"070d0765",	x"07320768",	
					x"07400774",	x"073b06c3",	x"213e5031",	x"06d0070e",	
					x"0708070f",	x"06d80715",	x"070a0714",	x"06ea0719",	
					x"06cf06fa",	x"06ce06fd",	x"06f006fe",	x"06bb0706",	
					x"06fa074f",	x"0711073a",	x"07310753",	x"070a072d",	
					x"0725072a",	x"07150742",	x"070f071c",	x"07060740",	
					x"073a073e",	x"0705074e",	x"0731075c",	x"07320774",	
					x"07450778",	x"07470766",	x"072d0738",	x"072d076a",	
					x"074e0762",	x"071f075c",	x"072a0796",	x"07370796",	
					x"0766078c",	x"07490776",	x"07480700",	x"213e6031",	
					x"06f90738",	x"06f80719",	x"06dc0728",	x"06e50713",	
					x"06df0706",	x"06df0709",	x"06f30705",	x"06dc0708",	
					x"06b80725",	x"06fc0734",	x"0707075d",	x"07340781",	
					x"0753077e",	x"07500773",	x"072b0779",	x"0744074f",	
					x"07430792",	x"07800789",	x"07760782",	x"0766079f",	
					x"07630797",	x"076f07a3",	x"07700793",	x"07600789",	
					x"07580780",	x"076207b1",	x"076107a1",	x"075707c3",	
					x"076707e3",	x"077907e4",	x"077e07e1",	x"077e0755",	
					x"213e7031",	x"072a0790",	x"07540760",	x"07380772",	
					x"0759076b",	x"07430745",	x"074b074a",	x"07360761",	
					x"07110734",	x"06e80799",	x"071d07a4",	x"075b07bf",	
					x"07a907d7",	x"079007f8",	x"079b07f1",	x"07ab07f7",	
					x"07b307be",	x"07b407f2",	x"07b107e2",	x"07bc07ff",	
					x"07f2081c",	x"07b70804",	x"07e80801",	x"07dd082d",	
					x"07e607d4",	x"07c20815",	x"07e707f0",	x"07eb07ee",	
					x"07f1083d",	x"07ea082b",	x"08060830",	x"07fb0826",	
					x"0810071d",	x"000a0004",	x"a3e84f0d",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"313f0031",	x"072b0732",	x"0743073e",	
					x"07360735",	x"07390738",	x"07140718",	x"070a0720",	
					x"070106fc",	x"06d806ac",	x"06d506de",	x"06ed06e2",	
					x"06ef06df",	x"074c0719",	x"07230734",	x"073d0744",	
					x"07450720",	x"072506f7",	x"07120717",	x"0746073d",	
					x"0757072d",	x"0752071b",	x"06fa070f",	x"06ff0733",	
					x"07210742",	x"07360701",	x"0726071a",	x"07320728",	
					x"073a0725",	x"072d0724",	x"0724074d",	x"071f0756",	
					x"072f0748",	x"073606ec",	x"313f1031",	x"071f0725",	
					x"074a0723",	x"07190706",	x"0714071e",	x"071606ea",	
					x"06f306ea",	x"06ee06bb",	x"06c406b0",	x"06a906d0",	
					x"06bb0703",	x"071306ff",	x"0717070c",	x"07160711",	
					x"0739072b",	x"07280727",	x"072906c8",	x"07080714",	
					x"07430727",	x"07260718",	x"073c0758",	x"07400719",	
					x"073b071a",	x"07120730",	x"07390702",	x"0718072d",	
					x"072b073c",	x"072e0720",	x"074a0720",	x"0709072d",	
					x"072d073e",	x"072d0749",	x"072306de",	x"313f2031",	
					x"070f06f7",	x"071906e6",	x"070f0703",	x"071e06f2",	
					x"06ef06df",	x"06db06e9",	x"06c506ae",	x"06ae0662",	
					x"069d06db",	x"06d806d1",	x"06f406e1",	x"06f406df",	
					x"06f00704",	x"07110708",	x"06f90712",	x"070d06e6",	
					x"07020737",	x"073906fe",	x"0708071d",	x"06f2071a",	
					x"07120721",	x"07230725",	x"07070708",	x"07180709",	
					x"06f80733",	x"070a0701",	x"07150719",	x"07290715",	
					x"06ed0711",	x"07150740",	x"07130740",	x"06fb06b3",	
					x"313f3031",	x"06bb06dc",	x"06d806e8",	x"06f1070e",	
					x"06fd0706",	x"06c106cf",	x"06bd06ea",	x"069906a7",	
					x"06b906b2",	x"06ad06c3",	x"068b06c4",	x"06c706ec",	
					x"06d30711",	x"06f70715",	x"07030718",	x"06f60723",	
					x"071806db",	x"06dd071f",	x"07130711",	x"06fa0718",	
					x"07190718",	x"07340727",	x"07230726",	x"0718071a",	
					x"0708071c",	x"06ea074c",	x"0721072f",	x"0704072d",	
					x"07010714",	x"07010722",	x"07100751",	x"07200746",	
					x"072006f7",	x"000a0004",	x"ce462591",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"31404031",	x"06c806f7",	x"06f60705",	
					x"06f90707",	x"0706070d",	x"06c906e7",	x"06f10704",	
					x"06af06d6",	x"06eb06d5",	x"06cc071f",	x"0709072e",	
					x"06f7072d",	x"0732073b",	x"06ec073f",	x"07200755",	
					x"07420758",	x"0732073f",	x"07370766",	x"07520770",	
					x"07650756",	x"07510766",	x"0757076f",	x"073a0752",	
					x"07420770",	x"075d073e",	x"0746076e",	x"0744077f",	
					x"075a0771",	x"07760780",	x"075d077c",	x"07690798",	
					x"07620799",	x"076e0722",	x"31405031",	x"072e0730",	
					x"074c074b",	x"072e076b",	x"075b0741",	x"070a077a",	
					x"072e074b",	x"0714071e",	x"07200727",	x"0722076c",	
					x"0749077e",	x"074e077b",	x"073f0779",	x"07390785",	
					x"07510787",	x"0767077e",	x"07590763",	x"0752078d",	
					x"07710793",	x"07620788",	x"075f07a0",	x"075e07a6",	
					x"076807ae",	x"076907bc",	x"07680793",	x"076b07c0",	
					x"077907b8",	x"076307d6",	x"077e07b5",	x"077f07c1",	
					x"077d07e0",	x"078c07ca",	x"07790732",	x"31406031",	
					x"0723074a",	x"07310756",	x"072f0762",	x"072d0747",	
					x"072f0751",	x"07460759",	x"070e0774",	x"0729074b",	
					x"07050778",	x"0739076b",	x"074a079d",	x"077507a2",	
					x"0762079f",	x"0778079a",	x"077f07b8",	x"077b0787",	
					x"077107ac",	x"078f07bb",	x"078f07be",	x"07b707d6",	
					x"079407c9",	x"079207ee",	x"079d07f3",	x"07b707c0",	
					x"079807e9",	x"07b307f4",	x"07b507ce",	x"079f080a",	
					x"079d080a",	x"0797081b",	x"07b0081b",	x"07ad074e",	
					x"31407031",	x"075107a6",	x"07700784",	x"076607c0",	
					x"0768079a",	x"076507a2",	x"0762078e",	x"0781077f",	
					x"075d0776",	x"075707c4",	x"07810800",	x"07af083b",	
					x"07c40816",	x"07cc0800",	x"07e90834",	x"07e2080a",	
					x"07f20828",	x"07f70832",	x"07fe0811",	x"08050841",	
					x"0815084b",	x"08220840",	x"0825086f",	x"083a0861",	
					x"0829082d",	x"08170865",	x"08230865",	x"082b0856",	
					x"0839085c",	x"082d0868",	x"0865087e",	x"08400854",	
					x"085a0680",	x"000a0004",	x"02186db5",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0241002e",	x"07400750",	x"07490746",	
					x"073a0726",	x"072f075a",	x"0754073d",	x"07480749",	
					x"07750758",	x"07700767",	x"078f079a",	x"07cc07af",	
					x"07890768",	x"07720776",	x"076e0780",	x"079b0784",	
					x"078f0775",	x"0797072c",	x"07840798",	x"079b078b",	
					x"0779078d",	x"07a50787",	x"075f0750",	x"0760077e",	
					x"07850769",	x"075e077a",	x"07ac0776",	x"07a6077e",	
					x"07780777",	x"07b30790",	x"078c0793",	x"07710792",	
					x"077e07a2",	x"07950725",	x"0241102e",	x"073c0726",	
					x"073e075d",	x"075d0706",	x"071e06fe",	x"0745073b",	
					x"0743075b",	x"075c075d",	x"076e0765",	x"07610772",	
					x"078a0796",	x"078a0759",	x"0772075d",	x"07540762",	
					x"078e077d",	x"0779077c",	x"07770757",	x"07560767",	
					x"07750761",	x"07510778",	x"07820771",	x"076e077f",	
					x"07aa0774",	x"078c0755",	x"0759076c",	x"078b075b",	
					x"07820787",	x"0795076d",	x"07800775",	x"077b077d",	
					x"07750765",	x"07840783",	x"0791071f",	x"0241202e",	
					x"0725072e",	x"072e0701",	x"070906f5",	x"072c0716",	
					x"0766073c",	x"0732072e",	x"0743072a",	x"0759073e",	
					x"0752076c",	x"076d075b",	x"07590742",	x"077c0751",	
					x"0764074f",	x"07560748",	x"0764073f",	x"07610745",	
					x"075b0754",	x"0763075d",	x"0765075f",	x"0766075e",	
					x"073d0747",	x"07320745",	x"07460755",	x"074a0743",	
					x"07750773",	x"07640753",	x"075a0733",	x"0751076f",	
					x"075d076d",	x"0758076d",	x"0757076c",	x"07500704",	
					x"0241302e",	x"06c40706",	x"070e071c",	x"072106f6",	
					x"06f40717",	x"070c0725",	x"07260748",	x"07390738",	
					x"07350712",	x"0718074b",	x"073e074d",	x"073a0744",	
					x"075c0734",	x"07340745",	x"0761073f",	x"0761075a",	
					x"074b072b",	x"072c0747",	x"073c074b",	x"074e0739",	
					x"073c075a",	x"0746073c",	x"0728074a",	x"073c0744",	
					x"074d073a",	x"074b077c",	x"07520777",	x"072e075f",	
					x"075c077c",	x"0758075c",	x"07420765",	x"07600781",	
					x"07640704",	x"000a0004",	x"3b724a87",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0242402e",	x"070b072d",	x"0708073a",	
					x"07150726",	x"070a072b",	x"071f071a",	x"0734072d",	
					x"07390735",	x"07440724",	x"073f0765",	x"07730761",	
					x"075a074f",	x"07520759",	x"074c0765",	x"075e075f",	
					x"07520771",	x"076c0759",	x"07610771",	x"07770784",	
					x"07780785",	x"07780782",	x"0794078b",	x"077f0790",	
					x"07840789",	x"07960764",	x"07a007aa",	x"07730787",	
					x"077f078d",	x"0796079d",	x"078307a8",	x"078007aa",	
					x"079107ad",	x"077e0750",	x"0242502e",	x"07360768",	
					x"0748078a",	x"075c0765",	x"0751076f",	x"074f076f",	
					x"078707a0",	x"078c07b1",	x"078b0782",	x"078a0797",	
					x"07840792",	x"079607a3",	x"07a807a6",	x"07a707aa",	
					x"079b0781",	x"079407c0",	x"079907a7",	x"079807c1",	
					x"07b607b1",	x"078007a7",	x"079d07a1",	x"078e07c8",	
					x"07a607bd",	x"078907c7",	x"07b107c0",	x"07b607d3",	
					x"079707c6",	x"079b07cf",	x"078807da",	x"07a307ca",	
					x"07aa07f7",	x"07b707f3",	x"07b4076b",	x"0242602e",	
					x"07300784",	x"0759075c",	x"075a0780",	x"075a078e",	
					x"07670771",	x"074b078b",	x"077307a8",	x"078707b0",	
					x"078e07c1",	x"07ba07be",	x"07ae07e1",	x"07b107e2",	
					x"07ab07cf",	x"07ba0805",	x"07bd07f3",	x"07db07cd",	
					x"07cb07eb",	x"07df07ee",	x"07d307e2",	x"07c507fd",	
					x"07c807ff",	x"07e707f4",	x"07f007e6",	x"07f507f2",	
					x"07d2081c",	x"07e807f2",	x"07ce0804",	x"07dc082e",	
					x"07d40825",	x"08060829",	x"07e40829",	x"07f2079c",	
					x"0242702e",	x"078307c3",	x"07a007b5",	x"07a007dd",	
					x"07c607dc",	x"07cc07bd",	x"07ce07f4",	x"081807fb",	
					x"07ee07ee",	x"07e2081e",	x"07f40831",	x"0813082e",	
					x"081e0841",	x"08180843",	x"08330835",	x"082d082d",	
					x"08440836",	x"0818085e",	x"08410874",	x"084e087d",	
					x"08520885",	x"0843084f",	x"08460880",	x"085f0864",	
					x"08570836",	x"0859086c",	x"088108b7",	x"086d0889",	
					x"086208c7",	x"088708bd",	x"088f08cd",	x"089308ac",	
					x"089d05d3",	x"000a0004",	x"664d82d4",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1243002e",	x"05e005d8",	x"05d705f5",	
					x"05fe05ea",	x"05fe05e8",	x"05f405e3",	x"05e20611",	
					x"062105df",	x"05ec05cf",	x"06050611",	x"0609061f",	
					x"06140628",	x"061e062d",	x"0653060c",	x"06160634",	
					x"063905ee",	x"061005d8",	x"0605061c",	x"063e0612",	
					x"06100621",	x"063c0629",	x"0628060a",	x"061d0617",	
					x"06090613",	x"06180605",	x"06060620",	x"06130632",	
					x"0628062e",	x"06140620",	x"0618061b",	x"06240621",	
					x"06010636",	x"060b05e1",	x"1243102e",	x"05ce05cc",	
					x"05d005c8",	x"05cc05df",	x"05e805e8",	x"05e705e4",	
					x"05e705f8",	x"05e705ee",	x"060105d0",	x"05ef0606",	
					x"060e0614",	x"0611060f",	x"061a0606",	x"061f0610",	
					x"06110619",	x"062705f7",	x"05fb05b8",	x"05fb05f7",	
					x"062805fb",	x"061205f9",	x"06070609",	x"061505fc",	
					x"061005fb",	x"060c060c",	x"061805f0",	x"05fd061a",	
					x"060d0617",	x"0613061a",	x"06160632",	x"061f062a",	
					x"06300627",	x"0623061b",	x"061b05b8",	x"1243202e",	
					x"05b105b2",	x"05d105cf",	x"05d505ca",	x"05df05ce",	
					x"05e405eb",	x"05fb05e5",	x"05f905e8",	x"05fc05d9",	
					x"060805dd",	x"05fe05e9",	x"06050600",	x"05f305f4",	
					x"05f105fc",	x"05fd05f8",	x"060505f4",	x"05f705ce",	
					x"05e205f1",	x"05fc05e6",	x"06010604",	x"061d05f7",	
					x"05e505ff",	x"05fb05fc",	x"05f605f8",	x"05fc05dc",	
					x"05df05e3",	x"06010616",	x"06000606",	x"05fb060d",	
					x"06000617",	x"0615060d",	x"05fa060d",	x"05f005c7",	
					x"1243302e",	x"05a605c7",	x"059d059d",	x"05aa05b2",	
					x"05bd05c9",	x"05e005c5",	x"05c405c6",	x"05c005e0",	
					x"05ca05a9",	x"05da05e7",	x"05db05e3",	x"05d405fa",	
					x"05ee05f8",	x"05f205f0",	x"05eb05f0",	x"05e605f4",	
					x"05dd05c0",	x"05d805fd",	x"05f405ee",	x"05f0060f",	
					x"05fd0606",	x"060405fc",	x"05fe060a",	x"05f405f5",	
					x"05eb05f4",	x"05f70605",	x"05f4060f",	x"06110615",	
					x"060b0617",	x"05fb0618",	x"06000616",	x"05fd061f",	
					x"060405d0",	x"000a0004",	x"cb019bd6",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1244402e",	x"05b005e0",	x"05c905db",	
					x"05c505e1",	x"05e20602",	x"05d405c1",	x"05e405da",	
					x"05de05da",	x"05eb05f1",	x"05ee05f0",	x"061c0607",	
					x"0619060f",	x"06150609",	x"05f9060a",	x"060305fe",	
					x"05f70605",	x"06070613",	x"05da0617",	x"0610061e",	
					x"062a0627",	x"062a061c",	x"0630062f",	x"062a061a",	
					x"06160625",	x"06280604",	x"06320634",	x"0631063e",	
					x"061f0635",	x"06470655",	x"0645063e",	x"0642065e",	
					x"06630652",	x"063505ff",	x"1244502e",	x"05e70612",	
					x"05f70602",	x"05f40623",	x"061a0626",	x"06220624",	
					x"05f20620",	x"06090648",	x"063a061a",	x"05fe063f",	
					x"062f0642",	x"062d0646",	x"0641065f",	x"06420650",	
					x"063f063d",	x"063c063c",	x"062a062b",	x"06170650",	
					x"0652064a",	x"06370650",	x"06430666",	x"06400659",	
					x"06420668",	x"0625066d",	x"064a0657",	x"06490644",	
					x"064e0682",	x"064f0675",	x"065c0688",	x"0651067a",	
					x"06620687",	x"0663068b",	x"06520635",	x"1244602e",	
					x"05eb0612",	x"05ee0611",	x"05ed0626",	x"061a062d",	
					x"06210640",	x"0603063d",	x"063a0649",	x"06260638",	
					x"06170659",	x"06460673",	x"064b0664",	x"06540667",	
					x"06510679",	x"06680665",	x"064b0661",	x"06580658",	
					x"065a066a",	x"0670067a",	x"06620685",	x"066906a4",	
					x"06970697",	x"06770692",	x"066d0698",	x"06800674",	
					x"0678069d",	x"067c069e",	x"068c06b4",	x"068506b2",	
					x"06760693",	x"067a06a6",	x"068a06bd",	x"06690650",	
					x"1244702e",	x"06160652",	x"06320640",	x"06240644",	
					x"06260687",	x"062e068e",	x"065e0679",	x"06650671",	
					x"0664068e",	x"065d06a5",	x"069606ca",	x"06a806ae",	
					x"069f06bd",	x"06bb06b7",	x"06bb06dd",	x"069a06b4",	
					x"06a10698",	x"06ad06cc",	x"06c906db",	x"06b506d3",	
					x"06b306e0",	x"06d406f3",	x"06ef06ed",	x"06c506dc",	
					x"06c306d0",	x"06dc06e3",	x"06cf06fc",	x"06f106f3",	
					x"06fd072d",	x"06fc0732",	x"0702071e",	x"0706070a",	
					x"06ed06d6",	x"000a0004",	x"f38cd10d",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2245002e",	x"06cd06ba",	x"06b306d2",	
					x"06f006e9",	x"06fa06ee",	x"06e106eb",	x"06ed06e6",	
					x"06fe070a",	x"06fa06fc",	x"06f806ee",	x"072f0709",	
					x"072506f2",	x"07290723",	x"070406f7",	x"07380707",	
					x"071906fd",	x"070806d5",	x"06df06e6",	x"06fb06f3",	
					x"06ee06d7",	x"0704070e",	x"0742071e",	x"072506d6",	
					x"06e006d9",	x"06e706e9",	x"06f206de",	x"06f50709",	
					x"06e806e7",	x"06f806f6",	x"06ee072b",	x"0717073f",	
					x"0707070e",	x"06f806a8",	x"2245102e",	x"06910690",	
					x"06a806c6",	x"06d206a5",	x"06bf06ad",	x"06da06cf",	
					x"06d006d0",	x"06e106d1",	x"06b506de",	x"06c906eb",	
					x"06fb06f6",	x"06fd06fe",	x"06fb06f0",	x"06fc06ed",	
					x"06eb06e7",	x"06f106e0",	x"06ee0691",	x"06c106d6",	
					x"06e306e9",	x"06fc06fa",	x"070a06fc",	x"070206f3",	
					x"06fb06e6",	x"06f206e6",	x"06ee06b6",	x"070606ec",	
					x"06fb06f6",	x"06fa06f9",	x"071a0719",	x"070b0710",	
					x"0711070b",	x"07090707",	x"0702068e",	x"2245202e",	
					x"068a0694",	x"069f06a4",	x"069e069d",	x"06b8069c",	
					x"06cb06b7",	x"06be06a7",	x"06ca06b7",	x"06d306b1",	
					x"06d406e5",	x"06fd06d6",	x"06fb06d6",	x"06e806d4",	
					x"06ea06c0",	x"06e306d5",	x"06df06d3",	x"06d706ad",	
					x"06c106b8",	x"06b606c3",	x"06c906df",	x"06d906ce",	
					x"06d606ea",	x"06fb06e5",	x"06e706da",	x"06cf06bc",	
					x"06cf06c6",	x"06ea06e4",	x"06ea06d1",	x"06dd06f6",	
					x"06c806d3",	x"06d906ed",	x"06ed06e8",	x"06d50667",	
					x"2245302e",	x"06580678",	x"0676068c",	x"06870699",	
					x"068f06a1",	x"069606ae",	x"06a4069c",	x"06c306ac",	
					x"06bc0691",	x"06ab06af",	x"06b806c3",	x"06d306ca",	
					x"06c806cf",	x"06cf06c2",	x"06c206ca",	x"06bc06c2",	
					x"06b50691",	x"068b06a7",	x"069f06b9",	x"06a506ab",	
					x"06c506bf",	x"06b806d1",	x"06dd06d2",	x"06d506da",	
					x"06d906c9",	x"06d006e5",	x"06c906cf",	x"06d606eb",	
					x"06d106ed",	x"06cd06f6",	x"06c806f5",	x"06d206f0",	
					x"06cc0672",	x"000a0004",	x"7b5f0a30",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2246402e",	x"06890693",	x"069c06aa",	
					x"06ca06a1",	x"06cb06ac",	x"06ae06bc",	x"06b606c0",	
					x"06db06ce",	x"06b706b7",	x"06c706dd",	x"06e906e0",	
					x"06e906cc",	x"06e106d0",	x"06dc06da",	x"06e706ec",	
					x"071006fa",	x"070506d5",	x"06ea06fb",	x"070006f5",	
					x"06f606f7",	x"06f20703",	x"06ed0703",	x"070a072e",	
					x"07130722",	x"06fc06e8",	x"0705071b",	x"070c0727",	
					x"07210727",	x"07150731",	x"071a072b",	x"07130727",	
					x"0710073f",	x"070f06ae",	x"2246502e",	x"069f06f4",	
					x"06d206da",	x"06e706ad",	x"06b706ce",	x"06e906f9",	
					x"06f806ec",	x"06f106fe",	x"070406f1",	x"06f8071c",	
					x"071f0732",	x"07000721",	x"07280716",	x"071c0713",	
					x"0715070f",	x"07010723",	x"070c06e0",	x"06f206f9",	
					x"070e071b",	x"07110721",	x"07140728",	x"070f0725",	
					x"07260741",	x"071e071e",	x"071d0733",	x"0726074d",	
					x"0735074e",	x"07190758",	x"0720075a",	x"0730076a",	
					x"073f076a",	x"0732075f",	x"073406c3",	x"2246602e",	
					x"06a506f8",	x"06b506e8",	x"06e906ed",	x"06f0070d",	
					x"06ea071d",	x"070c0722",	x"07110728",	x"0722071b",	
					x"07120755",	x"07510723",	x"072a0720",	x"07250759",	
					x"073c0753",	x"07440769",	x"07310750",	x"0743071f",	
					x"071f073a",	x"07520747",	x"07460766",	x"07530764",	
					x"076d0763",	x"07620771",	x"07640767",	x"0765076f",	
					x"07450775",	x"074c0793",	x"075507a6",	x"077907af",	
					x"07840797",	x"076f07a5",	x"077a07a4",	x"07790719",	
					x"2246702e",	x"070c0724",	x"070a0712",	x"0715071b",	
					x"07120755",	x"071f0724",	x"07340766",	x"07620748",	
					x"07440755",	x"076d0783",	x"0790078f",	x"07840785",	
					x"07a70790",	x"07970786",	x"078607cc",	x"07a30795",	
					x"07b80794",	x"078507bd",	x"07b407cf",	x"078d07eb",	
					x"08070808",	x"07bd07c6",	x"07c807ce",	x"07b107d4",	
					x"07c107d9",	x"07de07c6",	x"07c907f1",	x"07cf07ec",	
					x"07d807cd",	x"07da0821",	x"080b082b",	x"08040811",	
					x"080b06d9",	x"000a0004",	x"a59a3dc1",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3247002e",	x"06d606d4",	x"06fc06fe",	
					x"06c806ac",	x"06c206bc",	x"06d606f0",	x"0706070e",	
					x"07220703",	x"070006e6",	x"07170722",	x"07370725",	
					x"071806f1",	x"07360719",	x"07230703",	x"071b072b",	
					x"071906fa",	x"070e06e2",	x"070006fa",	x"07220704",	
					x"070f0712",	x"07120702",	x"06fe0711",	x"0724073b",	
					x"0734072e",	x"073906f5",	x"06ef0701",	x"070a0707",	
					x"07060708",	x"07170725",	x"0714070e",	x"07180728",	
					x"072a0706",	x"071e06dc",	x"3247102e",	x"06bf06af",	
					x"06b806c4",	x"06bc06c8",	x"06e206d4",	x"06d106da",	
					x"06d806f1",	x"06f206e0",	x"06ea06f2",	x"06fc06ff",	
					x"070a0713",	x"071f06ed",	x"06ec070b",	x"070e06c9",	
					x"06dd06e3",	x"06ea06eb",	x"06f306a6",	x"06de06d1",	
					x"06e406d2",	x"06bd06f1",	x"07020714",	x"070606ea",	
					x"06fb06f2",	x"06ff070f",	x"070206d5",	x"06ea06ee",	
					x"06f8070d",	x"06ef06db",	x"06ed070e",	x"070b070c",	
					x"07290726",	x"07360735",	x"073006da",	x"3247202e",	
					x"06d006a8",	x"06c6069f",	x"06ac06af",	x"06d906d4",	
					x"06de06d0",	x"070a06d5",	x"070a06de",	x"06fb06bc",	
					x"06f606f4",	x"071006f3",	x"070c06e3",	x"070706f2",	
					x"06fa06db",	x"06f606eb",	x"06e706d5",	x"06dc06b1",	
					x"06c106da",	x"06ea06db",	x"06c406d8",	x"06e206e4",	
					x"06c206f9",	x"06dc06f7",	x"06f206e7",	x"06df06d4",	
					x"06f706e0",	x"06e406e2",	x"06ef06e7",	x"06f606ff",	
					x"06ff06f5",	x"06e40702",	x"06ea06f0",	x"06df0690",	
					x"3247302e",	x"068d0684",	x"069b069e",	x"068a06a0",	
					x"06c106a9",	x"06ba06ac",	x"06b006ba",	x"06af06b1",	
					x"06bd06a1",	x"06d006cf",	x"06cb06b3",	x"06cb06dd",	
					x"06d906cd",	x"06cf06c1",	x"06ad06a3",	x"06a906bc",	
					x"06bc0696",	x"06bb06c5",	x"06b906b9",	x"06ba06c0",	
					x"06d706e6",	x"06c606ec",	x"06db06d7",	x"06d506e6",	
					x"06e306ba",	x"06c906de",	x"06d906ea",	x"06de06e0",	
					x"06d306f4",	x"06e006fc",	x"06df0700",	x"06e706ee",	
					x"06cd06b4",	x"000a0004",	x"c29d1170",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3248402e",	x"0685067e",	x"069006dc",	
					x"06ae06a3",	x"06b306b3",	x"06c006b6",	x"06ba06c2",	
					x"06e406bc",	x"06f506b1",	x"06e606d4",	x"06e506f5",	
					x"070906f6",	x"070706e7",	x"06d306fa",	x"06f606fb",	
					x"06ef06db",	x"06f406db",	x"06de06f9",	x"06f706f2",	
					x"07130702",	x"0728070b",	x"06f20708",	x"07080709",	
					x"0710071a",	x"071a0707",	x"0724070b",	x"07090706",	
					x"0712071b",	x"0725072d",	x"071e072c",	x"07140731",	
					x"07170722",	x"072806db",	x"3248502e",	x"06ba06d0",	
					x"06e206da",	x"06b906c9",	x"06c306e5",	x"06d206fc",	
					x"07170703",	x"072b0723",	x"07290705",	x"071b0719",	
					x"07110727",	x"0719073c",	x"0737072a",	x"071a073a",	
					x"071f070c",	x"07010704",	x"07190701",	x"0717072a",	
					x"0737071e",	x"070d073c",	x"07270738",	x"07150748",	
					x"072f0753",	x"073a0760",	x"07340721",	x"07220740",	
					x"07210750",	x"07250753",	x"07350775",	x"07580777",	
					x"07380761",	x"07380756",	x"071606cd",	x"3248602e",	
					x"06b406e4",	x"06f906dc",	x"06ac06f2",	x"06d006f6",	
					x"06d106f6",	x"0708071e",	x"072c072e",	x"071e0726",	
					x"070b0737",	x"07390753",	x"0739074b",	x"0740073b",	
					x"0723072d",	x"0725072d",	x"072b0740",	x"07350734",	
					x"0738075e",	x"07640762",	x"074a0757",	x"073a076a",	
					x"074e075f",	x"075d077a",	x"07520789",	x"0767074b",	
					x"07610761",	x"07600776",	x"07580783",	x"077e07ab",	
					x"078007b8",	x"07850797",	x"076e079b",	x"07720722",	
					x"3248702e",	x"072506f7",	x"06fc06fc",	x"06f70735",	
					x"072e0764",	x"074e074e",	x"073d0757",	x"07600748",	
					x"074e0765",	x"07590786",	x"07b107da",	x"07950792",	
					x"078207af",	x"079007a0",	x"079507c2",	x"07a807a9",	
					x"07b9077b",	x"07910791",	x"079b07b9",	x"07a707b9",	
					x"07c307e7",	x"07de07e7",	x"07dc07e3",	x"07dc07d7",	
					x"07f307cb",	x"07d007e0",	x"07e307e5",	x"07fd07ea",	
					x"080f0827",	x"08130834",	x"08150835",	x"083a0807",	
					x"080307b6",	x"000a0004",	x"e9564076",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0249002f",	x"07a607bf",	x"079507b8",	
					x"07a30791",	x"07960799",	x"0797078f",	x"077a07ad",	
					x"07a80785",	x"079f0726",	x"07530758",	x"075a0767",	
					x"07780736",	x"07540748",	x"07570762",	x"07900795",	
					x"079c076e",	x"07a30749",	x"0778078d",	x"079b0797",	
					x"07a8079a",	x"07b407a7",	x"078f077e",	x"07840790",	
					x"07790794",	x"077b0778",	x"0792077e",	x"07a9078e",	
					x"078a07a3",	x"07bf0772",	x"0777077f",	x"0764077e",	
					x"076c07a8",	x"077d0783",	x"0249102f",	x"07ab077e",	
					x"0790076d",	x"07820791",	x"07a80779",	x"07940757",	
					x"0773077a",	x"0778074c",	x"073f071f",	x"07240759",	
					x"07520758",	x"074f0719",	x"07420746",	x"073e0731",	
					x"073e0777",	x"0759074a",	x"075a0762",	x"074e0770",	
					x"07710774",	x"07710789",	x"07840795",	x"07aa075e",	
					x"078d07a2",	x"07bd0798",	x"0781077d",	x"07940777",	
					x"0777077f",	x"076e0792",	x"07810796",	x"07a207a2",	
					x"078f0786",	x"077f077f",	x"078a0757",	x"0249202f",	
					x"0769075b",	x"076a076c",	x"0771076c",	x"07980759",	
					x"07490762",	x"0765073f",	x"074d0768",	x"0785072a",	
					x"07390743",	x"075a0723",	x"072706fd",	x"07480723",	
					x"07390745",	x"076c0741",	x"07610742",	x"0769074b",	
					x"07630780",	x"076e0768",	x"075f076e",	x"076a0763",	
					x"0744076a",	x"07630770",	x"076e077c",	x"0769072b",	
					x"07570761",	x"076e0769",	x"0776076b",	x"07730777",	
					x"0775075b",	x"074e0769",	x"07730773",	x"075f0748",	
					x"0249302f",	x"074b076c",	x"077c075f",	x"075d0768",	
					x"073d0758",	x"0742074f",	x"0743074d",	x"074b0762",	
					x"0738072f",	x"070e072a",	x"072c0722",	x"070b071e",	
					x"071c0710",	x"07260743",	x"074c0742",	x"07510749",	
					x"07480740",	x"0748073c",	x"07500759",	x"07550756",	
					x"0758075c",	x"07600750",	x"0742075d",	x"074b0766",	
					x"07490742",	x"0742075a",	x"0754076a",	x"0741075c",	
					x"076f075f",	x"0748075d",	x"07430760",	x"0748078f",	
					x"075d0752",	x"000a0004",	x"41e05251",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"024a402f",	x"0745074c",	x"07260756",	
					x"073a0751",	x"074b0775",	x"074d0750",	x"074c077a",	
					x"0753073e",	x"074d0741",	x"073b0755",	x"07480747",	
					x"075c074d",	x"07520766",	x"074b0771",	x"0767077d",	
					x"076e076d",	x"07870777",	x"0771078b",	x"079207b0",	
					x"078a07a9",	x"07a60790",	x"07ae0776",	x"07790798",	
					x"07a70787",	x"078a076f",	x"078907ae",	x"079c079f",	
					x"07a0079c",	x"07a80799",	x"078607ab",	x"078d07b1",	
					x"078e07b0",	x"078f07a2",	x"024a502f",	x"077c07b2",	
					x"079d07b2",	x"07b607b9",	x"07b007b9",	x"0786079f",	
					x"077f079b",	x"078d079b",	x"07900793",	x"078f0789",	
					x"07800792",	x"07880763",	x"076f07ac",	x"079407af",	
					x"079707b1",	x"07a207ab",	x"079807b7",	x"079407c4",	
					x"07ad07b1",	x"077907a9",	x"079907c2",	x"07bb07d8",	
					x"07b507df",	x"07b107e0",	x"07b307cc",	x"07a307d4",	
					x"07aa07ea",	x"07ba07c9",	x"079c07ce",	x"078f07d9",	
					x"079f07ef",	x"07bf07eb",	x"07bb07bf",	x"024a602f",	
					x"079107d6",	x"07bb07b4",	x"078f07aa",	x"078c07ae",	
					x"078307c2",	x"079707cd",	x"079407b4",	x"079e07c0",	
					x"077107ca",	x"078907a2",	x"07500792",	x"078607d9",	
					x"076607d2",	x"07b407e1",	x"07aa07f3",	x"07bf07e1",	
					x"07bd0809",	x"080e080c",	x"07ee07e6",	x"07de080d",	
					x"07e20803",	x"07da0804",	x"07df07df",	x"07cb0810",	
					x"07e40835",	x"07ea0809",	x"07dd0816",	x"07ed0805",	
					x"07d1084b",	x"07fa084c",	x"07f60818",	x"07de07d5",	
					x"024a702f",	x"07bf07f4",	x"07d807ff",	x"07ad07d7",	
					x"07bb0803",	x"080207fc",	x"077707da",	x"07a007e8",	
					x"07c207e1",	x"0799080c",	x"07d507e7",	x"07a907e5",	
					x"07c4082b",	x"07e207f7",	x"07ec0839",	x"0810083a",	
					x"081e0855",	x"080e085b",	x"0856085a",	x"08160866",	
					x"084e0852",	x"085a0856",	x"0843089b",	x"0859086b",	
					x"0853086c",	x"086a0886",	x"0825088f",	x"08840871",	
					x"085f0899",	x"08600893",	x"086e08b7",	x"08780893",	
					x"088705f6",	x"000a0004",	x"67fa88b9",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"124b002f",	x"05fe0604",	x"0618060a",	
					x"062a05f4",	x"05eb05ea",	x"05e705e3",	x"05e505d5",	
					x"05ce05c0",	x"05d505b7",	x"05da05e2",	x"05fb0604",	
					x"06270649",	x"06280620",	x"06340607",	x"062e0613",	
					x"061f060d",	x"063905e4",	x"05ec062f",	x"06340603",	
					x"0621061b",	x"06320621",	x"06040610",	x"061b0638",	
					x"0627062a",	x"061e05f8",	x"060405ff",	x"060b0625",	
					x"060f0613",	x"062a062f",	x"0615063f",	x"062d0647",	
					x"06230639",	x"06230603",	x"124b102f",	x"05f005ea",	
					x"05e805ec",	x"05ef05df",	x"05d805d8",	x"05cc05ba",	
					x"05c305cb",	x"05cf05d1",	x"05d905c2",	x"05cd0600",	
					x"06080622",	x"06140620",	x"062a0624",	x"06190618",	
					x"06190620",	x"061505fb",	x"061105d7",	x"05ee0605",	
					x"06230600",	x"060d060f",	x"062505f8",	x"05fa05fb",	
					x"0607060b",	x"06060617",	x"05f805df",	x"05fb060f",	
					x"061d0608",	x"0619060f",	x"061f061e",	x"06200632",	
					x"0638063a",	x"062b0627",	x"062205c2",	x"124b202f",	
					x"05de05d0",	x"05ec05f5",	x"05cf05bb",	x"05dd05ce",	
					x"05d105d2",	x"05e705ac",	x"05c605ae",	x"05bc05ad",	
					x"05dd05d6",	x"05db05de",	x"05ea0601",	x"05f105e7",	
					x"05fe05f4",	x"060605fc",	x"05fe05f7",	x"05df05cf",	
					x"05df05ed",	x"05e905f2",	x"06000601",	x"06140602",	
					x"05f70605",	x"05fb05f0",	x"05f40617",	x"060005e6",	
					x"05fa0607",	x"06040614",	x"0605060d",	x"05f3061e",	
					x"05fb060e",	x"060f060a",	x"05f40614",	x"061505c4",	
					x"124b302f",	x"05a805d4",	x"05d405e2",	x"05c005c7",	
					x"05a105dd",	x"05c305bb",	x"05a405c7",	x"05cc05c6",	
					x"05af05b0",	x"05d105e1",	x"05e705e0",	x"05e005e8",	
					x"05e405f9",	x"05e705f8",	x"05ea0604",	x"05ec05ed",	
					x"05eb05ce",	x"05dc05fb",	x"06070619",	x"06080618",	
					x"06040614",	x"05fd060d",	x"0610061b",	x"060a05ff",	
					x"05f705f0",	x"0605061f",	x"06000616",	x"05ee0622",	
					x"060d0629",	x"05fe0631",	x"061a0633",	x"06140637",	
					x"061e05f4",	x"000a0004",	x"caca9d57",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"124c402f",	x"05e105ea",	x"05cf05f4",	
					x"05ef05e6",	x"05bf05e1",	x"05a405e5",	x"05ca05d2",	
					x"05d005d1",	x"05d305e0",	x"05a20601",	x"06030618",	
					x"061e0626",	x"0609061a",	x"0606061d",	x"061e0623",	
					x"06150626",	x"061c061e",	x"06110635",	x"062a062e",	
					x"06130645",	x"06440642",	x"063c0655",	x"064b064d",	
					x"063d0648",	x"06370619",	x"06270663",	x"064f0655",	
					x"0623066d",	x"064e0675",	x"064c0669",	x"064f066d",	
					x"065b0677",	x"064b05f3",	x"124c502f",	x"05df062a",	
					x"05f50630",	x"05fe0620",	x"06000621",	x"0603061c",	
					x"0608062b",	x"05d90633",	x"05f50616",	x"05ff0650",	
					x"06260652",	x"0629064e",	x"065b065e",	x"062e064f",	
					x"06300658",	x"063d0661",	x"06260630",	x"06230663",	
					x"065a0673",	x"06530675",	x"06570675",	x"06570697",	
					x"065b0680",	x"064a0671",	x"06420659",	x"063e0697",	
					x"06600699",	x"06520692",	x"06590696",	x"06520680",	
					x"065806a1",	x"0663068c",	x"0650060c",	x"124c602f",	
					x"05e4064c",	x"06000623",	x"05fa062c",	x"06190634",	
					x"05f00635",	x"05ec0651",	x"05fe061f",	x"05f70653",	
					x"061c065c",	x"0638065c",	x"06430666",	x"06580668",	
					x"06520695",	x"0669068e",	x"06700695",	x"067f0664",	
					x"064d068f",	x"06820684",	x"066906a8",	x"0678069f",	
					x"068706ac",	x"069606a2",	x"069706b9",	x"066d0687",	
					x"068a06ae",	x"068506b2",	x"068006cb",	x"069d06ba",	
					x"068806ba",	x"068206bc",	x"068806bf",	x"06750636",	
					x"124c702f",	x"0611065e",	x"063d0656",	x"06340683",	
					x"062d069b",	x"060f067d",	x"063e0681",	x"06350650",	
					x"06360687",	x"0627068a",	x"065806cd",	x"067e06e9",	
					x"069e06d7",	x"06a306d8",	x"06bc06c0",	x"06bc06e0",	
					x"06a206a6",	x"069106f8",	x"06e60707",	x"06b006fe",	
					x"06e60708",	x"06b90712",	x"06e606f3",	x"06d106f0",	
					x"06c506ba",	x"06cc06ff",	x"06d306f2",	x"06df0707",	
					x"07070733",	x"06f5073b",	x"06f40711",	x"0704072f",	
					x"06fd06df",	x"000a0004",	x"f359d962",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"224d002f",	x"06e106db",	x"06b706e7",	
					x"06c306bd",	x"06cd06d3",	x"06c106be",	x"06d806d9",	
					x"06cd06ea",	x"06db06b4",	x"06bc06c9",	x"06ea0703",	
					x"071006f3",	x"07200707",	x"07080702",	x"07220708",	
					x"071106fe",	x"071d06d3",	x"06f706e0",	x"06ea0707",	
					x"07010715",	x"07280704",	x"07060719",	x"07110729",	
					x"071406ed",	x"06fc06db",	x"070106f4",	x"07130722",	
					x"070c0717",	x"07070716",	x"06ef0717",	x"0706071f",	
					x"06f90710",	x"070a06cf",	x"224d102f",	x"06e206c9",	
					x"06ee06be",	x"06b506c0",	x"06e8069c",	x"069306c2",	
					x"06bf06bd",	x"06d606c4",	x"06c706ad",	x"06c006e5",	
					x"06e606f1",	x"070406f1",	x"070206f7",	x"071606fe",	
					x"06fb06ca",	x"06d806d9",	x"06df06c6",	x"06c506cf",	
					x"06d906d1",	x"06dc06e5",	x"06f30700",	x"06ef0716",	
					x"071806df",	x"070006e9",	x"070206d8",	x"070d0707",	
					x"070e0700",	x"06f406fb",	x"07130725",	x"070c0715",	
					x"071a0701",	x"0708071b",	x"07070688",	x"224d202f",	
					x"06a90689",	x"06a306be",	x"06c706bd",	x"06c3069a",	
					x"06a90691",	x"06af06b4",	x"06c606b1",	x"06b706a2",	
					x"06c006bf",	x"06e806e1",	x"070606e2",	x"06e006d2",	
					x"06e006d6",	x"06ce06c9",	x"06dc06da",	x"06eb06ca",	
					x"06e806e6",	x"06db06dd",	x"06d606ef",	x"06e206cb",	
					x"06df06d5",	x"06d006f8",	x"06e006f2",	x"06db06be",	
					x"06d606e6",	x"06e406e7",	x"06e606e8",	x"06e506e5",	
					x"06d1070d",	x"06f006fa",	x"06e606ee",	x"06dd0698",	
					x"224d302f",	x"06690686",	x"066006a6",	x"06730693",	
					x"067c0697",	x"0681069b",	x"06a106ae",	x"06a3068e",	
					x"067f0664",	x"068106bf",	x"06ca06c6",	x"06be06c2",	
					x"06c206cf",	x"06cd06d1",	x"06c206de",	x"06bc06cc",	
					x"06c3069d",	x"06c306bb",	x"06cb06e3",	x"06c806db",	
					x"06e106e5",	x"06ca06ef",	x"06d406e7",	x"06df06f8",	
					x"06e406ce",	x"06bb06f5",	x"06c406e7",	x"06d106ee",	
					x"06d106f0",	x"06d00713",	x"06ca070b",	x"06e50707",	
					x"06ea06aa",	x"000a0004",	x"7b3a0d65",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"224e402f",	x"068406ba",	x"06ac06bf",	
					x"069706a7",	x"06a206e5",	x"069a06c7",	x"06a006c0",	
					x"06b606ec",	x"06b306ac",	x"06bd06ef",	x"06d106fe",	
					x"071006ec",	x"06fd06f3",	x"06e006f4",	x"06f6071f",	
					x"07010704",	x"06fe06e7",	x"06d90702",	x"06f2072c",	
					x"070f071c",	x"070a0716",	x"07090725",	x"07080721",	
					x"071d0724",	x"071e0710",	x"07210739",	x"0728074a",	
					x"0725074b",	x"0741074e",	x"0727073e",	x"07270739",	
					x"070f074f",	x"072f06d9",	x"224e502f",	x"06b1070a",	
					x"06db0724",	x"06c906ef",	x"06e40700",	x"06d80711",	
					x"06e606fa",	x"06cb0714",	x"06e506fc",	x"06fd072c",	
					x"0708074b",	x"07250738",	x"071d0720",	x"071b0750",	
					x"0741073f",	x"07010754",	x"07220724",	x"07230740",	
					x"07180745",	x"07290764",	x"07340748",	x"070b0761",	
					x"07350753",	x"071d0753",	x"071d074e",	x"0722076c",	
					x"072a0771",	x"072f0769",	x"073a076e",	x"073f077d",	
					x"073b076e",	x"07390779",	x"073b06f3",	x"224e602f",	
					x"06c1070d",	x"06e20710",	x"0706070b",	x"06d206f9",	
					x"06a906fb",	x"06bc0708",	x"06ec074e",	x"06fb0725",	
					x"06e70757",	x"07190766",	x"0752076a",	x"0753076d",	
					x"073b0785",	x"076a07ae",	x"0749077f",	x"0732074d",	
					x"0723077f",	x"07510779",	x"075b0782",	x"075607a6",	
					x"076e07a5",	x"07620785",	x"075b0782",	x"075d076e",	
					x"075d07a2",	x"075b07a3",	x"075307a8",	x"076807b1",	
					x"076c07b1",	x"076d07b4",	x"076f07a8",	x"075f075f",	
					x"224e702f",	x"06fa0742",	x"06f40708",	x"06f70726",	
					x"0718073a",	x"07170743",	x"0711073d",	x"070a0737",	
					x"071e0772",	x"074107ab",	x"0785077b",	x"077107b3",	
					x"077a07b3",	x"079d07c6",	x"07ad07cd",	x"077a07c4",	
					x"0791077e",	x"076b07de",	x"07ce07fc",	x"07bb0802",	
					x"07e5081c",	x"07ce0817",	x"07ee0808",	x"07c70804",	
					x"07b80801",	x"07f00812",	x"07ed07fe",	x"07e207f9",	
					x"07e10808",	x"08060828",	x"07d50820",	x"07fe0811",	
					x"080c06fa",	x"000a0004",	x"a5704bdc",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"324f002f",	x"06f706d9",	x"06f506dd",	
					x"06e606b8",	x"06b206c6",	x"06b606d0",	x"06d00708",	
					x"06e00706",	x"070d06ba",	x"06d20720",	x"07070724",	
					x"07270721",	x"073006d8",	x"06e30703",	x"0718070f",	
					x"07470700",	x"073506ed",	x"070906ea",	x"07070750",	
					x"072e0724",	x"072e0721",	x"070e0710",	x"071d0720",	
					x"0722070a",	x"071c0712",	x"0720071d",	x"072a0739",	
					x"0719070e",	x"06f50703",	x"070f0711",	x"07100734",	
					x"07270719",	x"070e06b7",	x"324f102f",	x"06cd06b8",	
					x"06d206bd",	x"06d306ac",	x"06c406bf",	x"06c106c9",	
					x"06d706e0",	x"06e606df",	x"06d906b7",	x"06df0719",	
					x"071d070e",	x"070406f0",	x"06f10707",	x"070206f9",	
					x"071d070e",	x"070406ff",	x"070306db",	x"070006e3",	
					x"0702070b",	x"072a06f8",	x"070606f7",	x"06f906f6",	
					x"073306f4",	x"071906eb",	x"06fa06cd",	x"06e806f9",	
					x"07040710",	x"07040712",	x"071a071d",	x"07040713",	
					x"07170717",	x"0728072f",	x"072706ab",	x"324f202f",	
					x"06bc06aa",	x"06bd06b1",	x"069d06b7",	x"06c006c6",	
					x"06da06c7",	x"070006d3",	x"06ef06c7",	x"06e206b3",	
					x"06eb06d1",	x"071406e7",	x"070206f0",	x"070406d8",	
					x"06e106ec",	x"06f206ce",	x"06db0700",	x"06e806c3",	
					x"06dc06e7",	x"06e706fc",	x"06f006f8",	x"06f006dd",	
					x"06d606ee",	x"06fd06fe",	x"06f50705",	x"06ee06d5",	
					x"06fb0709",	x"06f706fd",	x"06e80708",	x"06f906e5",	
					x"06e40702",	x"06fe0704",	x"06e80720",	x"06ec0684",	
					x"324f302f",	x"0675068b",	x"067f068d",	x"06750680",	
					x"069c06a1",	x"068506a6",	x"06a306ab",	x"068806b5",	
					x"06cd0696",	x"06b406d5",	x"06c706c3",	x"06c906d8",	
					x"06c006df",	x"06e006dd",	x"06d606d3",	x"06da06c5",	
					x"06ce06a6",	x"06df06e2",	x"06cd06eb",	x"06cc06e8",	
					x"06f306fe",	x"06de0704",	x"06f206fb",	x"06f706f8",	
					x"06e806f4",	x"070a071a",	x"070e0701",	x"06e606fd",	
					x"06e80712",	x"06f10701",	x"06db0702",	x"06e7070f",	
					x"06eb06cb",	x"000a0004",	x"c45314a8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3250402f",	x"068906c1",	x"06aa06b5",	
					x"068a06be",	x"06c106a6",	x"069f06be",	x"06c706c7",	
					x"06c606ca",	x"06f006cc",	x"06dd0707",	x"06eb070c",	
					x"06fb0717",	x"07070704",	x"06fa070e",	x"06fb071f",	
					x"07130720",	x"071106f1",	x"06fe072a",	x"07090720",	
					x"073a0731",	x"071e072e",	x"0719072c",	x"071f0728",	
					x"071e074b",	x"071a0724",	x"073d0775",	x"07300745",	
					x"072c074e",	x"07300734",	x"07150752",	x"071b0763",	
					x"07410767",	x"071906e5",	x"3250502f",	x"06e80704",	
					x"06d706fa",	x"06c306fe",	x"06c40714",	x"06cd0711",	
					x"07050704",	x"06f30733",	x"072a070f",	x"07230736",	
					x"07200755",	x"07500751",	x"07480740",	x"072a0745",	
					x"072f0745",	x"07390748",	x"071a0728",	x"0725076a",	
					x"0744076d",	x"07380753",	x"07280752",	x"072b0766",	
					x"073d0778",	x"073907a6",	x"07470752",	x"0741079b",	
					x"074d076f",	x"074e0776",	x"074b0781",	x"075407a3",	
					x"075f077e",	x"076007ad",	x"074d06fd",	x"3250602f",	
					x"06db072c",	x"06e8071f",	x"06d206e9",	x"06dc072c",	
					x"06ea0723",	x"06ff071b",	x"06f0072d",	x"071d0726",	
					x"07110776",	x"07370789",	x"073b0778",	x"0745078f",	
					x"072b0780",	x"0759077e",	x"0751077e",	x"0784076c",	
					x"07460782",	x"0760078f",	x"076b0794",	x"07560794",	
					x"07570784",	x"077e07a3",	x"076c07b3",	x"07710781",	
					x"07740792",	x"077e07b5",	x"078107ba",	x"078a07b1",	
					x"077b07e3",	x"079007e1",	x"078f07e2",	x"0771073a",	
					x"3250702f",	x"07050738",	x"07160736",	x"07010745",	
					x"07030786",	x"07170752",	x"0726074f",	x"07160756",	
					x"073b0759",	x"073e07af",	x"077807b5",	x"077b07c2",	
					x"07b007b2",	x"079907cf",	x"077e07d4",	x"07a307e4",	
					x"077e07b5",	x"078a07ea",	x"07b007ec",	x"07a40807",	
					x"07e30832",	x"07cf07fd",	x"07f20802",	x"07f2081c",	
					x"07dc07e6",	x"07ea0820",	x"07fa0818",	x"080a0817",	
					x"07e1083d",	x"08080839",	x"07fe0847",	x"07fd0827",	
					x"07ef0603",	x"000a0004",	x"ed435225",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"02510030",	x"06f608c0",	x"06c907ca",	
					x"07b20503",	x"03e7062f",	x"05ae079c",	x"08c80692",	
					x"0839071d",	x"076e0482",	x"07180883",	x"0861052f",	
					x"08cc045f",	x"08950855",	x"07d70894",	x"08fc0691",	
					x"07b608a1",	x"0504059d",	x"06d50592",	x"03a40583",	
					x"067d0882",	x"07070575",	x"04d70704",	x"07e2070f",	
					x"089206c8",	x"07b5056a",	x"0518082b",	x"061a072d",	
					x"060c0846",	x"0943068d",	x"064f06b2",	x"05cc07e9",	
					x"05fa02fc",	x"063f06e0",	x"02511030",	x"08a9069b",	
					x"06af0732",	x"06c607fd",	x"08c205d9",	x"05a3053c",	
					x"07ba0477",	x"082308cc",	x"06e30325",	x"04d805e1",	
					x"0584061f",	x"086505bf",	x"074d0687",	x"074807dd",	
					x"06ca0433",	x"056605b1",	x"05b5085b",	x"080e062f",	
					x"06760652",	x"06d1075f",	x"062806e9",	x"076403cd",	
					x"05de05a8",	x"06df0747",	x"05bf04df",	x"0705048d",	
					x"064d06b8",	x"068d0651",	x"08490818",	x"05ee0679",	
					x"0650075f",	x"082b0861",	x"04ec07dc",	x"02512030",	
					x"048007be",	x"07dc07cb",	x"07ea07dd",	x"082e07d4",	
					x"080a07cd",	x"07d407c2",	x"07d407be",	x"08150805",	
					x"081307fe",	x"081e07c8",	x"07aa07a9",	x"07b007a7",	
					x"07ae0790",	x"07b507c2",	x"076e07c3",	x"07f007e8",	
					x"058d07a7",	x"079007ad",	x"076f07c1",	x"07c80755",	
					x"077406b5",	x"076407a8",	x"07870712",	x"075e07cf",	
					x"06d50555",	x"0730070f",	x"07d9059f",	x"078a07f2",	
					x"082507e0",	x"07dd07bf",	x"07e30822",	x"080007d7",	
					x"02513030",	x"07c007aa",	x"07de07ff",	x"07ea07d2",	
					x"07c107d2",	x"07cc07c8",	x"07aa07de",	x"07e307d6",	
					x"07df07ec",	x"07d8079c",	x"07b507ae",	x"07aa078d",	
					x"07c207a3",	x"07980783",	x"07a607a5",	x"07c607bc",	
					x"07ba07f2",	x"079c0746",	x"079307b8",	x"079207ba",	
					x"07800775",	x"07ae0777",	x"076b0786",	x"0797078d",	
					x"07c307d7",	x"07ac07bd",	x"079007c6",	x"07c707d5",	
					x"07e207e0",	x"07e20803",	x"07e707fa",	x"07d20800",	
					x"07e907bf",	x"000a0004",	x"2d732c0c",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"02524030",	x"07a607de",	x"07d607ee",	
					x"07e607e5",	x"07e307f8",	x"081307e9",	x"07ed07f6",	
					x"07f407f7",	x"080a0824",	x"082b07ce",	x"07e207c2",	
					x"07d907a2",	x"07c907c7",	x"07d507dd",	x"07d207c9",	
					x"07c907f4",	x"08070804",	x"07e407dd",	x"07e107e2",	
					x"07d507ee",	x"07b807e9",	x"07f507d7",	x"07ca07e6",	
					x"07dd07e0",	x"07f50819",	x"08010804",	x"07ff07fe",	
					x"07fd07f5",	x"0812082a",	x"081f0842",	x"08310836",	
					x"0827085e",	x"083c0828",	x"02525030",	x"07f3083c",	
					x"083a0863",	x"08560862",	x"08520840",	x"083f083d",	
					x"085a085b",	x"085e0844",	x"085f0858",	x"0834082f",	
					x"08170823",	x"081e0804",	x"080b0801",	x"08070806",	
					x"0801080b",	x"08030835",	x"08330824",	x"0808081e",	
					x"080f07ea",	x"07c707e9",	x"07e307fc",	x"07e40805",	
					x"07d6081b",	x"07ef085c",	x"08390855",	x"083e0854",	
					x"0828084b",	x"0823084c",	x"0800086f",	x"083f0883",	
					x"084f089c",	x"085f0897",	x"08680844",	x"02526030",	
					x"0808084e",	x"08660864",	x"08600868",	x"085c0870",	
					x"085f0871",	x"086b0879",	x"0864085e",	x"085e087c",	
					x"08400845",	x"0856083d",	x"08400838",	x"082f0843",	
					x"07f30828",	x"08190844",	x"081e0856",	x"08520885",	
					x"08650843",	x"084a0852",	x"083a0848",	x"083d085c",	
					x"08140839",	x"08430859",	x"0849086a",	x"082c08a4",	
					x"087108af",	x"0856087b",	x"08460891",	x"085508b5",	
					x"087e08be",	x"08af08d1",	x"089108d7",	x"088f08c7",	
					x"02527030",	x"087108bc",	x"08c408f5",	x"08ce08b6",	
					x"08da08cf",	x"08e008dd",	x"08e208ce",	x"08da08b5",	
					x"08cf08ff",	x"08dd08c0",	x"08d708aa",	x"08aa08b8",	
					x"08a908bb",	x"089f08b3",	x"08b608ac",	x"08ad08b0",	
					x"08dc08da",	x"08bb087c",	x"089608d4",	x"089f0908",	
					x"08c408c6",	x"08a008bc",	x"08b80913",	x"08dc08bd",	
					x"08cc0913",	x"091408fc",	x"08e8093d",	x"091a0933",	
					x"08f20958",	x"09170966",	x"094a0961",	x"09560953",	
					x"093f05c2",	x"000a0004",	x"b45bcd49",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"12530030",	x"05cd05ce",	x"05dd05e0",	
					x"060805f0",	x"05fb05fc",	x"05ec05ec",	x"05f505ff",	
					x"06110611",	x"061505cc",	x"060b060c",	x"0618061c",	
					x"0610061a",	x"062905f9",	x"061a05f9",	x"060605fb",	
					x"061405ff",	x"060905de",	x"05e90602",	x"06210606",	
					x"060d0605",	x"06030609",	x"06060607",	x"06100609",	
					x"05f4060a",	x"062205d8",	x"05e6060f",	x"0608061c",	
					x"062d061e",	x"0621063c",	x"061c0639",	x"06380632",	
					x"05fa0636",	x"062005db",	x"12531030",	x"05f305cd",	
					x"05da05ce",	x"05d105dc",	x"05d105ee",	x"05fd05ee",	
					x"05f105fa",	x"06160613",	x"062405df",	x"05ef05f8",	
					x"0613060d",	x"060c060f",	x"06120617",	x"061c060e",	
					x"061c0605",	x"060d0601",	x"05e205d1",	x"05ed05e0",	
					x"060405fa",	x"06120607",	x"062205f7",	x"060905f8",	
					x"05fb0619",	x"06170611",	x"060605e2",	x"0604062f",	
					x"062a061c",	x"062d062a",	x"0632061e",	x"060b0629",	
					x"06360628",	x"06160621",	x"062f05c1",	x"12532030",	
					x"05c305bd",	x"05d005da",	x"05c605d2",	x"05d305ca",	
					x"05bc05bd",	x"060505fb",	x"06050607",	x"060505e7",	
					x"060105f1",	x"060b05fa",	x"061a0605",	x"05fc05f4",	
					x"060605e3",	x"05e405e9",	x"05eb05dd",	x"05ec05b7",	
					x"05ce05ef",	x"05f105ff",	x"05fb060b",	x"060f0607",	
					x"05f90604",	x"060d05fe",	x"06020609",	x"05ff05da",	
					x"05b605ff",	x"05f7060d",	x"05fd060c",	x"06020619",	
					x"06080616",	x"06160605",	x"05fb0619",	x"05f905b4",	
					x"12533030",	x"05eb05ba",	x"05a305c4",	x"05c205d4",	
					x"05d305e6",	x"05dd05e3",	x"05f205cb",	x"05e005f1",	
					x"05ef05b4",	x"05e405de",	x"05df05f8",	x"05ff05f4",	
					x"05e805f2",	x"05ec05e2",	x"05f00600",	x"05e705d6",	
					x"05b805ac",	x"05c605ec",	x"05fe05f9",	x"05f90607",	
					x"05fe0612",	x"060005f2",	x"05fe05f8",	x"05d205fe",	
					x"05fc05f1",	x"05dc0617",	x"06050605",	x"06000610",	
					x"05f80619",	x"0601062f",	x"0614062f",	x"0612062b",	
					x"05fb05db",	x"000a0004",	x"cb7e9c4a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"12544030",	x"05d505e0",	x"05e10602",	
					x"05de05ec",	x"05df0607",	x"05dc0603",	x"05ff05e6",	
					x"05e605f5",	x"05fc0600",	x"05fd05ff",	x"061a0609",	
					x"06210604",	x"06090605",	x"05fe060a",	x"06190605",	
					x"060805fe",	x"060f05f6",	x"060f061d",	x"060a0635",	
					x"063a0643",	x"0641064f",	x"0635063c",	x"062f062f",	
					x"0623062b",	x"0624061e",	x"061c0627",	x"0629064f",	
					x"063d064f",	x"065a0659",	x"06490655",	x"0640064d",	
					x"065c066f",	x"065b0608",	x"12545030",	x"05f5061b",	
					x"06000636",	x"05eb0621",	x"0617062f",	x"062a0638",	
					x"06230636",	x"063b0635",	x"064b0639",	x"061d064a",	
					x"064a0656",	x"064c064a",	x"064a065f",	x"064a065a",	
					x"06530656",	x"06340644",	x"0632063d",	x"062d064f",	
					x"06480657",	x"06550652",	x"0649065e",	x"0655066a",	
					x"0657067b",	x"063a0677",	x"06510659",	x"063f0659",	
					x"065d0688",	x"06550671",	x"065c0698",	x"06630689",	
					x"06850688",	x"065d0678",	x"0655063f",	x"12546030",	
					x"0608062b",	x"06140632",	x"0608062e",	x"060e0642",	
					x"06360647",	x"062d0665",	x"06480662",	x"0651065e",	
					x"064f066b",	x"06570679",	x"06510664",	x"0668067a",	
					x"066a067b",	x"066b0664",	x"065c0686",	x"066b0671",	
					x"064b067e",	x"06670676",	x"06710694",	x"0688069e",	
					x"068306aa",	x"06720694",	x"068006a0",	x"06910687",	
					x"06800687",	x"067d068f",	x"067e06ba",	x"069606b5",	
					x"068e06b9",	x"068c06ae",	x"069506b6",	x"0683067d",	
					x"12547030",	x"0642068c",	x"065b0679",	x"0633067f",	
					x"067b06b3",	x"067606bb",	x"068b06bb",	x"068e06b3",	
					x"06a106a1",	x"068406cd",	x"06c806d5",	x"06be06d1",	
					x"06cc06c8",	x"06bc06d9",	x"06d206d2",	x"06bb06bf",	
					x"06cc06a5",	x"06c406f6",	x"06db0704",	x"06dc06f9",	
					x"06e206f1",	x"06f30707",	x"06f806f7",	x"070106f9",	
					x"06f606c7",	x"06d906fd",	x"06eb070c",	x"06e8070d",	
					x"0718073f",	x"07150745",	x"07360744",	x"07070720",	
					x"071606c5",	x"000a0004",	x"fd22d911",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"22550030",	x"06ec06af",	x"06c706cb",	
					x"06c306cb",	x"06de06d9",	x"06e306e1",	x"06ff0727",	
					x"073706f2",	x"06f006c5",	x"06c9070a",	x"071c070c",	
					x"06f806e2",	x"071d071e",	x"070306d9",	x"06fe06ef",	
					x"070f06fe",	x"06ff06b5",	x"06e306dc",	x"070406f5",	
					x"06ee06df",	x"06f806e6",	x"07150719",	x"07160708",	
					x"07020705",	x"06ef06c6",	x"06da06ec",	x"070706f5",	
					x"06f806ee",	x"06fb072e",	x"07080721",	x"0702070d",	
					x"0707072b",	x"07030699",	x"22551030",	x"06ab06aa",	
					x"06c006dc",	x"06db06ae",	x"06ca06a3",	x"06c906b6",	
					x"06d906e8",	x"070606f1",	x"06f106a9",	x"06ec06f9",	
					x"06f306f5",	x"06ee06ed",	x"06fa06f4",	x"06f106f5",	
					x"06fd06d1",	x"06e006ca",	x"06ec06c1",	x"06bc06e4",	
					x"06f606f4",	x"071106ee",	x"070306d2",	x"06ec0716",	
					x"0706070c",	x"070506e7",	x"06e006a6",	x"06e506f6",	
					x"06eb06db",	x"06e006fe",	x"06f2071a",	x"0714072f",	
					x"072406f5",	x"06fe0723",	x"071506be",	x"22552030",	
					x"06c906a8",	x"06a7067d",	x"06b506a2",	x"06bb06a8",	
					x"06b106a1",	x"06d606cc",	x"06ce06c2",	x"06d4067f",	
					x"06d306d9",	x"06f106d2",	x"06e906d0",	x"06df06c8",	
					x"06df06d4",	x"06f806c4",	x"06bb06c8",	x"06dc0671",	
					x"06b706bd",	x"06ba06cb",	x"06c806cd",	x"06cb06c1",	
					x"069606fa",	x"06ec06f4",	x"06dc06ef",	x"06d006c5",	
					x"06c706d7",	x"06dd06d4",	x"06da06e2",	x"06ea06e0",	
					x"06db06e5",	x"06d206f8",	x"06e406f2",	x"06dd066b",	
					x"22553030",	x"068c069b",	x"069f0698",	x"06870693",	
					x"0690069e",	x"069c06b2",	x"06b406b3",	x"06ce0688",	
					x"06ac0676",	x"06b706b7",	x"06d206d2",	x"06c806d0",	
					x"06b806d5",	x"06c206ca",	x"06bc06c6",	x"06b206ac",	
					x"06b00691",	x"06a806a5",	x"06c106c2",	x"06af06c4",	
					x"06ca06cb",	x"06b706d9",	x"06e506d6",	x"06db06eb",	
					x"06cc06b7",	x"06c206fd",	x"06cf06ce",	x"06cf06fa",	
					x"06ec06f9",	x"06d6070d",	x"06be06fc",	x"06ce06f9",	
					x"06df0685",	x"000a0004",	x"7be00abd",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"22564030",	x"06950678",	x"068a06c8",	
					x"06b906b4",	x"06ba06c4",	x"06b306b4",	x"06a206c1",	
					x"06d906c9",	x"06d306d2",	x"06d906e6",	x"06e006e3",	
					x"06f406de",	x"06ed06f5",	x"06f206cd",	x"06f006f7",	
					x"06ef06ee",	x"06f506e9",	x"06f706fe",	x"071f06ff",	
					x"07150703",	x"070206f5",	x"06fb0703",	x"06f50715",	
					x"07090709",	x"07050703",	x"07060712",	x"07080717",	
					x"0711071e",	x"0719072e",	x"07120722",	x"07170737",	
					x"071b073f",	x"073406d7",	x"22565030",	x"06e506fa",	
					x"06f306ea",	x"06fc06de",	x"06bf070c",	x"06dc06e6",	
					x"06e506fb",	x"06fd0715",	x"070e0709",	x"0713071a",	
					x"072c0736",	x"072e0720",	x"071f0711",	x"0720070b",	
					x"07140711",	x"07130710",	x"06f806ee",	x"06dc0720",	
					x"0720072e",	x"07110746",	x"073c0737",	x"070a0739",	
					x"0724074e",	x"072c0731",	x"071e0731",	x"07290764",	
					x"07330756",	x"072e0751",	x"073c077f",	x"073d0772",	
					x"0741075e",	x"0744075f",	x"074a06e4",	x"22566030",	
					x"06d806fc",	x"06f10703",	x"06ea0707",	x"06f10737",	
					x"070a0714",	x"0706071e",	x"07130723",	x"072e0739",	
					x"07330756",	x"07500760",	x"07520733",	x"07430750",	
					x"07510754",	x"07480767",	x"07350766",	x"07410747",	
					x"07370741",	x"07570777",	x"076f0784",	x"076e076e",	
					x"07630781",	x"075b078c",	x"077a0788",	x"077b0771",	
					x"076d0783",	x"076a078f",	x"075d0796",	x"077a07b8",	
					x"077907aa",	x"077b07b1",	x"078f07b7",	x"077d0721",	
					x"22567030",	x"07380765",	x"0732072d",	x"07280770",	
					x"075a0788",	x"077007a5",	x"079b0791",	x"078a077e",	
					x"07830778",	x"077807b7",	x"07d307d3",	x"07cd07b3",	
					x"07b807ba",	x"07c307b1",	x"07a907d9",	x"07c507bc",	
					x"07bf07b1",	x"07b607ca",	x"07d907fe",	x"07db07f7",	
					x"07ff080c",	x"07e407fb",	x"080307f4",	x"07e707e1",	
					x"07cf07e0",	x"07ea07f4",	x"07f30821",	x"07f3080e",	
					x"08010840",	x"0809083b",	x"0844084b",	x"081f0819",	
					x"083206ce",	x"000a0004",	x"aef446ef",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"32570030",	x"06f806b2",	x"06d006de",	
					x"06d006b1",	x"06c706b2",	x"06d206a9",	x"06cd06f1",	
					x"06e806f0",	x"071006e6",	x"071406d8",	x"070b0702",	
					x"070f06f9",	x"071b06f1",	x"07070720",	x"070d06f8",	
					x"07040710",	x"072a06c1",	x"06df06ee",	x"07080710",	
					x"06fb06f3",	x"070606f7",	x"06fc0703",	x"06e40709",	
					x"0707070e",	x"06fc06e6",	x"06ed06f6",	x"07180709",	
					x"06f606eb",	x"06d206fd",	x"07070707",	x"070b0735",	
					x"072806f7",	x"06fa06b0",	x"32571030",	x"06ae067a",	
					x"06a406a2",	x"06be067f",	x"06cb06be",	x"06dc06b3",	
					x"06d406eb",	x"06dd06f9",	x"06f506c3",	x"06d706fb",	
					x"070506e1",	x"06e806bf",	x"06dc0734",	x"070506d3",	
					x"06ef06ee",	x"06e806d9",	x"06ee06ba",	x"06ef06d5",	
					x"06f706dc",	x"06e006e5",	x"06e706e7",	x"06f706d2",	
					x"06f906e2",	x"06fa06ef",	x"06f606e1",	x"06d406f1",	
					x"06eb06f4",	x"06e006f2",	x"06f906fc",	x"06fb071a",	
					x"07210728",	x"072c071a",	x"071206b8",	x"32572030",	
					x"06df069d",	x"06b206a3",	x"06b106ad",	x"06b506aa",	
					x"06c206ca",	x"06fc06c4",	x"06dd06e0",	x"070606a1",	
					x"06fa06c8",	x"070106d8",	x"070d06f4",	x"070806ed",	
					x"06f906d8",	x"06ee06cb",	x"06c706cb",	x"06cd06af",	
					x"06c106ed",	x"06f406d7",	x"06d006da",	x"06d506e1",	
					x"06ca06db",	x"06e106fc",	x"070706ff",	x"06f3069c",	
					x"06bb06c0",	x"06d206db",	x"06d006e3",	x"06e406e9",	
					x"06e706f1",	x"06f00724",	x"07060703",	x"06ef068b",	
					x"32573030",	x"06a50684",	x"06950690",	x"06970698",	
					x"069a069d",	x"069206be",	x"068806cb",	x"06dc06bc",	
					x"06cf06a2",	x"06e406da",	x"06c806c0",	x"06c806ce",	
					x"06c806cc",	x"06ce06d0",	x"06ce06ad",	x"06b706a8",	
					x"06ac0693",	x"06bb06af",	x"06b106d3",	x"06b906bf",	
					x"06ce06c6",	x"06c806d8",	x"06d606e2",	x"06e906ea",	
					x"06d906b7",	x"06b306d0",	x"06ca06d2",	x"06d406dc",	
					x"06e206fe",	x"06f00706",	x"06ea0708",	x"06ef06f6",	
					x"06d506ad",	x"000a0004",	x"be9c0c06",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"32584030",	x"06ad06a1",	x"069e06b9",	
					x"068c06a0",	x"06a6069c",	x"06a306b4",	x"06cd06c0",	
					x"06c706c2",	x"06ee06bc",	x"06dd06ec",	x"06f206e1",	
					x"070606e5",	x"06ec06e9",	x"06ee0709",	x"06f506f0",	
					x"070106f6",	x"06fb06c6",	x"06e306e7",	x"06f10700",	
					x"07240701",	x"0734070c",	x"070606fe",	x"06f606f8",	
					x"0705070c",	x"071306fb",	x"071c071a",	x"07170725",	
					x"071d0728",	x"07270734",	x"071b073c",	x"07340744",	
					x"07340743",	x"072906c0",	x"32585030",	x"06df06e4",	
					x"070006e2",	x"06aa06e0",	x"06fa06f1",	x"06f406fb",	
					x"071806f7",	x"07290721",	x"07300718",	x"072d072e",	
					x"0720072c",	x"07280728",	x"07250711",	x"071c0702",	
					x"070f0718",	x"0714072e",	x"071306ff",	x"07170730",	
					x"0736072f",	x"0736072d",	x"07170747",	x"07100750",	
					x"07360769",	x"07490758",	x"073e0735",	x"07230745",	
					x"073e073b",	x"073f0754",	x"073e077a",	x"07500784",	
					x"07530772",	x"074d0769",	x"07350704",	x"32586030",	
					x"0702070b",	x"06d706f2",	x"06e506f4",	x"06d00728",	
					x"070e0725",	x"072c071d",	x"072d0731",	x"07330740",	
					x"07320748",	x"072e0761",	x"073d074b",	x"075a075a",	
					x"073c0750",	x"07480748",	x"074f076d",	x"074d0733",	
					x"07470758",	x"07570763",	x"074f075c",	x"07470776",	
					x"07630774",	x"07810796",	x"0767077c",	x"076d0753",	
					x"07590795",	x"0768078b",	x"076107a7",	x"078207a1",	
					x"077807b0",	x"079507ae",	x"079607ac",	x"07790741",	
					x"32587030",	x"07550736",	x"07320764",	x"0750076e",	
					x"076a0783",	x"074b0769",	x"07390798",	x"078707a1",	
					x"07970782",	x"076007cc",	x"07cc07dc",	x"07d007a4",	
					x"07c107cf",	x"07b807c4",	x"07bb07e6",	x"07c007e9",	
					x"07e607a0",	x"07b507e0",	x"07bc07df",	x"07df07d1",	
					x"07d407fb",	x"07ee07ef",	x"07ea07f0",	x"07ff0807",	
					x"080707e2",	x"07e20808",	x"08070808",	x"07fb0807",	
					x"0813083b",	x"08170836",	x"0818083c",	x"082b0817",	
					x"08140761",	x"000a0004",	x"f13e47e0",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"02590031",	x"0796079a",	x"078b0789",	
					x"07780767",	x"076307a0",	x"077e077c",	x"0780077c",	
					x"07780740",	x"07540721",	x"07440732",	x"07350740",	
					x"072b073f",	x"0758072f",	x"07320744",	x"07600779",	
					x"0789073a",	x"0777075c",	x"077b077d",	x"079a078e",	
					x"07780784",	x"07a1079e",	x"0769077e",	x"0785077d",	
					x"0776076c",	x"076a074f",	x"0760076e",	x"07720773",	
					x"0757075a",	x"07770764",	x"076a0761",	x"07420760",	
					x"07660767",	x"075d071a",	x"02591031",	x"07630748",	
					x"07630737",	x"07750749",	x"07620763",	x"075e074f",	
					x"075f0748",	x"073c072e",	x"0739070c",	x"0708070e",	
					x"070d0720",	x"070e0709",	x"07260755",	x"073a0725",	
					x"07370740",	x"07250748",	x"07530759",	x"07400744",	
					x"07610778",	x"076c0778",	x"07780760",	x"07780760",	
					x"07790778",	x"07750751",	x"0752071d",	x"07430741",	
					x"07550740",	x"07560747",	x"0755077d",	x"07770791",	
					x"07700778",	x"077b0768",	x"0774072f",	x"02592031",	
					x"0744074b",	x"074c0744",	x"075f0753",	x"074f074a",	
					x"0742072d",	x"0723070d",	x"070f072d",	x"073406f8",	
					x"0723072d",	x"07200709",	x"07070706",	x"07420705",	
					x"072c0731",	x"07240726",	x"07400736",	x"07540732",	
					x"07420785",	x"076c075b",	x"07610752",	x"075f0759",	
					x"07320750",	x"0739074d",	x"0741075a",	x"0745071d",	
					x"073c0764",	x"07450750",	x"07600742",	x"07450743",	
					x"074b074c",	x"07410759",	x"07410743",	x"07370710",	
					x"02593031",	x"070b0722",	x"0723072d",	x"0723072d",	
					x"0711071c",	x"07150734",	x"07220728",	x"070506f8",	
					x"06f106f2",	x"06d90705",	x"072006f8",	x"06d3070e",	
					x"070506ed",	x"07070707",	x"0727072c",	x"073c0725",	
					x"0723072a",	x"072a072f",	x"073a0747",	x"0757074c",	
					x"073d0754",	x"07510739",	x"07310740",	x"073b0744",	
					x"07240710",	x"07030747",	x"0741074e",	x"0729074e",	
					x"07560760",	x"0743074d",	x"072f0744",	x"073b075a",	
					x"07350715",	x"000a0004",	x"31534240",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"025a4031",	x"074e0742",	x"07350739",	
					x"07340745",	x"07450740",	x"07260732",	x"072d0748",	
					x"072c072f",	x"072e0703",	x"070a0727",	x"07050716",	
					x"070f072b",	x"071f0735",	x"072a0761",	x"075f075c",	
					x"07640769",	x"07760768",	x"07660783",	x"078c078e",	
					x"07800787",	x"07770782",	x"07920774",	x"07930791",	
					x"07800779",	x"076a076e",	x"077307ac",	x"0784079c",	
					x"0783077b",	x"079d0791",	x"0793079b",	x"077c0793",	
					x"07720796",	x"076f076c",	x"025a5031",	x"07760789",	
					x"07670767",	x"076d0780",	x"076a0788",	x"07540773",	
					x"07670768",	x"075c0782",	x"07540757",	x"07620767",	
					x"0755076b",	x"07640770",	x"0779077e",	x"07780794",	
					x"078e079b",	x"0781079c",	x"078a07a2",	x"078707b5",	
					x"079607c5",	x"0768079f",	x"079807ca",	x"07bd07d3",	
					x"07ab07c6",	x"079a07c4",	x"07a707bc",	x"077d07d7",	
					x"078f07c8",	x"079207d3",	x"078407d6",	x"078c07ea",	
					x"07ab07ec",	x"07b707e6",	x"07ac077f",	x"025a6031",	
					x"0775079b",	x"0778079e",	x"0791079a",	x"07770799",	
					x"0779079f",	x"078207a2",	x"0781078b",	x"0750075f",	
					x"07460783",	x"07730788",	x"075d0794",	x"078e07b2",	
					x"077d07c5",	x"07ad07d5",	x"07b207df",	x"07bd07cb",	
					x"07bc0805",	x"07f207f3",	x"07e007f6",	x"07ee0816",	
					x"07e507fa",	x"07d407f7",	x"07e7081e",	x"07f207e3",	
					x"07b5081c",	x"08030815",	x"07da07f7",	x"07d20807",	
					x"07de081f",	x"08000823",	x"07e60816",	x"07d607ee",	
					x"025a7031",	x"07f807fc",	x"07cd0811",	x"07d50809",	
					x"07e6081d",	x"08000814",	x"07f40821",	x"07b307fe",	
					x"07bd07e2",	x"07b207c5",	x"07d607d3",	x"07c507ea",	
					x"07e6083a",	x"07ce080c",	x"07ef082c",	x"0823084c",	
					x"08420861",	x"081b0868",	x"08540866",	x"08500875",	
					x"085e088e",	x"0876085b",	x"0867088d",	x"0883087c",	
					x"0878087c",	x"08780884",	x"0875089d",	x"087f089b",	
					x"089b08d4",	x"086a08b4",	x"088e08be",	x"089e089c",	
					x"089c05f8",	x"000a0004",	x"64578220",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"125b0031",	x"05fc05e7",	x"05fb05fd",	
					x"05f705c0",	x"05d705d5",	x"05d305b9",	x"05df05e6",	
					x"05db05aa",	x"05cd05c8",	x"05e205df",	x"05f50604",	
					x"05ff05fe",	x"060e0627",	x"06360619",	x"06330614",	
					x"0641061b",	x"0616060b",	x"06070612",	x"062b060d",	
					x"06110604",	x"06100605",	x"06120601",	x"06050624",	
					x"0603060c",	x"0616060a",	x"05fc0600",	x"060d0620",	
					x"061d0613",	x"06340613",	x"0607063b",	x"06290644",	
					x"0622062a",	x"061605df",	x"125b1031",	x"05eb05e8",	
					x"05e705dc",	x"05df05ea",	x"05dd05be",	x"05ab05ca",	
					x"05b005a0",	x"05a705d4",	x"05e905be",	x"05cf05e1",	
					x"05fb0607",	x"05f20614",	x"06080631",	x"061305fe",	
					x"05fe05fa",	x"060d05f9",	x"061505cf",	x"05ee05f3",	
					x"05fd0603",	x"06160609",	x"061105fd",	x"060a05fd",	
					x"060d0601",	x"060a05f7",	x"061005d1",	x"05f8060d",	
					x"05fb0603",	x"06210617",	x"061c0604",	x"060c061c",	
					x"06200622",	x"061f0614",	x"060b05b8",	x"125b2031",	
					x"05ea05cd",	x"05e405e0",	x"05cc05c0",	x"05c805c9",	
					x"05ae05b6",	x"05d305ab",	x"05d105c7",	x"05dd05bb",	
					x"05d005c1",	x"05db05e7",	x"05f005fc",	x"05e405ec",	
					x"05ef0616",	x"060b05f2",	x"05ef05ec",	x"05fe05dd",	
					x"05dc05e6",	x"05ea05e3",	x"05fa0606",	x"06090600",	
					x"05e80603",	x"060105ff",	x"060105fc",	x"060005be",	
					x"05e605f4",	x"05f805fb",	x"05e80603",	x"06070614",	
					x"06030611",	x"06110607",	x"06010613",	x"05f605d3",	
					x"125b3031",	x"05be05a8",	x"05ae05ad",	x"05a705de",	
					x"05d405d6",	x"05ba05c0",	x"05a105b9",	x"05aa05c2",	
					x"059c05ac",	x"05c205e5",	x"05dc05e8",	x"05dd05f5",	
					x"05fa05fd",	x"05f205fa",	x"05f10600",	x"05f105f8",	
					x"05f305cb",	x"05b30609",	x"05f30610",	x"05f8060e",	
					x"05f80615",	x"060f060d",	x"0602060d",	x"05f60621",	
					x"05e705eb",	x"05e30624",	x"05fc0615",	x"05f40627",	
					x"06140623",	x"05ff0627",	x"060f0631",	x"0611062f",	
					x"05ff05de",	x"000a0004",	x"c76a99c1",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"125c4031",	x"05d605f7",	x"05db05fe",	
					x"05e705e9",	x"05d405e5",	x"05c705e3",	x"05cd05e5",	
					x"05cf05d8",	x"05d505ee",	x"05c905f2",	x"05eb060d",	
					x"06140637",	x"06270621",	x"06140626",	x"062b062e",	
					x"06100639",	x"061e0606",	x"06190638",	x"062d063a",	
					x"06350645",	x"06390650",	x"063e0649",	x"063a063f",	
					x"06320633",	x"0632062d",	x"06270652",	x"06450659",	
					x"0639064b",	x"06440650",	x"0644065a",	x"06530659",	
					x"06580662",	x"06410616",	x"125c5031",	x"05fe0640",	
					x"06180625",	x"05d70624",	x"0602060b",	x"06090623",	
					x"06150629",	x"060a0630",	x"0603061f",	x"061d065d",	
					x"06460666",	x"06480648",	x"064c0658",	x"063a065f",	
					x"065a0655",	x"061f0654",	x"06380650",	x"063a0669",	
					x"06520673",	x"063b0673",	x"064e0671",	x"0651068f",	
					x"065a0691",	x"064e0678",	x"06570671",	x"06570680",	
					x"065d069b",	x"06480683",	x"065e06b4",	x"065906ac",	
					x"066d0699",	x"06780683",	x"06680633",	x"125c6031",	
					x"062a062e",	x"06160642",	x"06180636",	x"06230642",	
					x"06250647",	x"06260634",	x"061f0641",	x"060f063d",	
					x"06150663",	x"061d0666",	x"06510681",	x"06620685",	
					x"065e068f",	x"06700697",	x"067d0688",	x"06880673",	
					x"06610690",	x"068f0681",	x"066e06a1",	x"068706a4",	
					x"069306b6",	x"068206a3",	x"068806b0",	x"0691068d",	
					x"067a06ab",	x"067b06b6",	x"069306cf",	x"069906c6",	
					x"068b06c8",	x"069d06c8",	x"069706b4",	x"067e0691",	
					x"125c7031",	x"0659068b",	x"06590687",	x"062d0675",	
					x"0648069e",	x"064b0697",	x"0640068c",	x"066106a6",	
					x"06680683",	x"066406e5",	x"068f06e3",	x"06a806e5",	
					x"06cf06e3",	x"069a06f3",	x"06e806f0",	x"06e106ee",	
					x"06c106c1",	x"06c1070b",	x"06d5071a",	x"06de070d",	
					x"06e30700",	x"06ef0721",	x"07010720",	x"06fe0714",	
					x"06ed06f9",	x"06f1071b",	x"07140729",	x"07090724",	
					x"071d0739",	x"07180754",	x"070e073e",	x"071b073c",	
					x"071206c8",	x"000a0004",	x"fb3fde0d",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"225d0031",	x"070506e2",	x"06c406c8",	
					x"06a806b2",	x"06b206b5",	x"06ac06c1",	x"06de06ed",	
					x"06e906d1",	x"06db06b8",	x"06c506dc",	x"06ff06e4",	
					x"06fd06ea",	x"071e070b",	x"070906f4",	x"07210716",	
					x"072506d9",	x"06ed06df",	x"070606de",	x"06f206f2",	
					x"06ed06f5",	x"06fc0712",	x"070a06f3",	x"070706eb",	
					x"070006d8",	x"06f506e3",	x"06f0071f",	x"071206f2",	
					x"06dc06ea",	x"06fe072c",	x"06ef070b",	x"07080730",	
					x"06d506e1",	x"06c90696",	x"225d1031",	x"06bc06b5",	
					x"06d106dd",	x"06d606b8",	x"06bb069a",	x"06a106d3",	
					x"06bf06be",	x"069206c5",	x"06c606c4",	x"06ce06d0",	
					x"06f6070d",	x"06f606f4",	x"06ed06ee",	x"06ec06e6",	
					x"06ee06ca",	x"06eb06d3",	x"06ca0696",	x"06ce06cf",	
					x"06d706e6",	x"06f806e4",	x"06ed06e2",	x"06e406f3",	
					x"06eb06e4",	x"06e706cd",	x"06e806b0",	x"06ef06d7",	
					x"06e8070a",	x"071206e5",	x"06fd0717",	x"06f0070d",	
					x"070406fe",	x"070106ea",	x"070e0691",	x"225d2031",	
					x"06c806b0",	x"06a706bb",	x"06d306a3",	x"06be06a0",	
					x"0696067d",	x"0686068f",	x"06980693",	x"06ad0689",	
					x"06b406d2",	x"06e706cd",	x"06f106df",	x"06d306b6",	
					x"06c706cf",	x"06fe06db",	x"06d506d0",	x"06d706c8",	
					x"06d406ce",	x"06cb06d5",	x"06e206e5",	x"06e106db",	
					x"06e306f8",	x"06e706e0",	x"06d406e3",	x"06ec06bb",	
					x"06ac06e0",	x"06dc06d8",	x"06d706ec",	x"06f406ed",	
					x"06da06fb",	x"06e506fa",	x"06eb06f3",	x"06e50694",	
					x"225d3031",	x"068a06b6",	x"066c06a1",	x"06690681",	
					x"06840690",	x"066b06c8",	x"068e06a1",	x"069706ab",	
					x"06ae0680",	x"0687068e",	x"06b006d2",	x"06d406ab",	
					x"06af06b3",	x"06b606e1",	x"06ba06dc",	x"06c906c4",	
					x"06c706ae",	x"06b206a7",	x"06b906df",	x"06c806ef",	
					x"06e0070e",	x"06c706e3",	x"06cf06d0",	x"06c306dc",	
					x"06c706e5",	x"06c406f2",	x"06c006dd",	x"06db06e9",	
					x"06d40705",	x"06dd0712",	x"06db0711",	x"06e906fb",	
					x"06da06d5",	x"000a0004",	x"781f0a72",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"225e4031",	x"069b06a7",	x"068906a6",	
					x"068706a4",	x"06a006dd",	x"069206cd",	x"06aa06c9",	
					x"06d806bf",	x"06af06a5",	x"06d006fe",	x"06d70704",	
					x"06e906ee",	x"06d006ff",	x"06f30711",	x"07070714",	
					x"07030709",	x"0711070d",	x"06f10711",	x"07130718",	
					x"071e0710",	x"06fd071e",	x"070b0723",	x"0721072a",	
					x"071d0724",	x"07010718",	x"07130730",	x"07240739",	
					x"0710073c",	x"07220751",	x"0731074e",	x"07300750",	
					x"0714074e",	x"071706f6",	x"225e5031",	x"06ce070c",	
					x"06f106ff",	x"06ea06e0",	x"06d106fb",	x"06ef0720",	
					x"06fe0709",	x"06fa0724",	x"07100700",	x"06d90720",	
					x"06fc0746",	x"07290741",	x"071c072d",	x"0729073d",	
					x"07290744",	x"071e0752",	x"07190730",	x"071d0747",	
					x"07270756",	x"073e074f",	x"07330746",	x"072e0760",	
					x"0733075b",	x"072c0756",	x"073a075d",	x"06f80772",	
					x"0738077b",	x"07350770",	x"07400772",	x"0745077d",	
					x"07370768",	x"07400771",	x"074106f5",	x"225e6031",	
					x"06eb074d",	x"06dd06f8",	x"06d2070b",	x"06dd0723",	
					x"0706071c",	x"06fa0728",	x"0706072d",	x"071c0745",	
					x"07130757",	x"0745076d",	x"0753075c",	x"0753076e",	
					x"0727078e",	x"076207a2",	x"07570794",	x"07640767",	
					x"074f0782",	x"078a0783",	x"075e0795",	x"075c0795",	
					x"076b0796",	x"075e07a0",	x"07730791",	x"07590785",	
					x"076907a0",	x"076407b1",	x"076b07cb",	x"078507c1",	
					x"078707c3",	x"077607b8",	x"078307a7",	x"078c0733",	
					x"225e7031",	x"073d075d",	x"07480765",	x"07400736",	
					x"07330797",	x"07410781",	x"072f075b",	x"07480761",	
					x"0761078e",	x"077c07cd",	x"079807bb",	x"07be07ec",	
					x"07c807f5",	x"07d40803",	x"07d307ff",	x"07b207df",	
					x"07c007ad",	x"07ae0812",	x"07e90831",	x"07e307fb",	
					x"07fd0841",	x"07dc081f",	x"07ec0809",	x"08010829",	
					x"07e407e9",	x"07d30834",	x"08190825",	x"081b0824",	
					x"081e083e",	x"081a085e",	x"0833084b",	x"08310835",	
					x"082806da",	x"000a0004",	x"aef3521a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"325f0031",	x"06e006b8",	x"06b806c0",	
					x"06c006b8",	x"06bc06b4",	x"06b306b1",	x"06b106cd",	
					x"06ca0709",	x"06d206cc",	x"06eb06e4",	x"06eb070d",	
					x"06fd06fa",	x"06fa0720",	x"071d06f5",	x"0719070b",	
					x"071f072d",	x"071806a2",	x"06d506da",	x"06f10709",	
					x"07100710",	x"07210704",	x"06f60715",	x"072806fe",	
					x"070d06ef",	x"071d06fe",	x"06fc0730",	x"0738072e",	
					x"0700071c",	x"07110702",	x"06ee06ef",	x"06f90726",	
					x"070b0703",	x"06f706ab",	x"325f1031",	x"06b906b0",	
					x"06c106bb",	x"06d206ae",	x"06f106ab",	x"06a306aa",	
					x"06a806b3",	x"06d706c2",	x"06d606a1",	x"06eb06eb",	
					x"06eb06e2",	x"06f006e7",	x"06f506f8",	x"06ef06e6",	
					x"070b06e5",	x"06e7070e",	x"06eb069f",	x"06d106bf",	
					x"06e306ed",	x"06e506ec",	x"070d06e4",	x"06e506e4",	
					x"07030702",	x"071606e6",	x"06f106b6",	x"07110702",	
					x"06eb071d",	x"0700071c",	x"06f606f8",	x"06eb0702",	
					x"06ee0707",	x"0714070d",	x"070c06b5",	x"325f2031",	
					x"06c206a7",	x"06a006a5",	x"069906ae",	x"06bd069f",	
					x"06cd06b6",	x"06d906c7",	x"06d006e0",	x"06e9069d",	
					x"06d206d5",	x"06f506e4",	x"070806cd",	x"06e606c3",	
					x"06da06d7",	x"06ed06bf",	x"06db06ea",	x"06ea06b0",	
					x"06b606d9",	x"06cb06f5",	x"06d406f6",	x"06e606df",	
					x"06bb06eb",	x"06fb06ec",	x"06e306ed",	x"06da06e0",	
					x"06e206ed",	x"06e306e9",	x"06d606eb",	x"070606f3",	
					x"06cb06eb",	x"06b806f8",	x"06e7070c",	x"06d20681",	
					x"325f3031",	x"068e069a",	x"06ab06b2",	x"068e0683",	
					x"0682068e",	x"068406c0",	x"069906c0",	x"06ac06ad",	
					x"06b60682",	x"06b506e2",	x"06ce06ba",	x"06c206c7",	
					x"06cc06cf",	x"06da06da",	x"06d906e1",	x"06dc06d9",	
					x"06dd06b5",	x"06c506cf",	x"06ba06e2",	x"06c906e0",	
					x"06fe06f0",	x"06fe06e9",	x"06e606f9",	x"06eb06e7",	
					x"06e406e2",	x"06d806fd",	x"06e706ed",	x"06e806f2",	
					x"06f10715",	x"06f10719",	x"06ee0718",	x"06e006fb",	
					x"06db06d5",	x"000a0004",	x"bdb50ea7",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"32604031",	x"06b506c5",	x"06a906a7",	
					x"06b206c1",	x"06b206a9",	x"06af06c3",	x"06d006c6",	
					x"06c406cf",	x"06e006a4",	x"06c606f3",	x"06df06fd",	
					x"070a070d",	x"070c070c",	x"06e2070e",	x"06ea070d",	
					x"06f50703",	x"070106fd",	x"06ff0718",	x"07140729",	
					x"073f072d",	x"0714073a",	x"07210739",	x"07240739",	
					x"07230737",	x"071b0714",	x"07230739",	x"072a073d",	
					x"072a072f",	x"072f0724",	x"07050726",	x"07160759",	
					x"07230760",	x"072006f4",	x"32605031",	x"06fb0701",	
					x"06e50708",	x"06d70703",	x"06f50739",	x"06ec0718",	
					x"07020717",	x"06fe072c",	x"07120721",	x"0720073c",	
					x"072b0743",	x"07450751",	x"07430748",	x"07390756",	
					x"0725074d",	x"07380740",	x"072d0727",	x"071d0737",	
					x"07400755",	x"071f075a",	x"07350766",	x"0716077e",	
					x"074e0783",	x"07400781",	x"07380762",	x"07320796",	
					x"07570771",	x"07430768",	x"0741077a",	x"07520799",	
					x"07590795",	x"075a077c",	x"074c06ea",	x"32606031",	
					x"06ed0736",	x"06f00713",	x"06d60729",	x"07030731",	
					x"06e2073f",	x"07200733",	x"071a073b",	x"07310732",	
					x"0715075a",	x"0729076f",	x"07610799",	x"076c0797",	
					x"074c076c",	x"07590777",	x"075c0784",	x"0767076c",	
					x"076d0783",	x"07790799",	x"077d079a",	x"076d07b0",	
					x"077707a2",	x"078f07be",	x"077d07ac",	x"077a078c",	
					x"0792079c",	x"079907dc",	x"079507bc",	x"079107ac",	
					x"077e07bb",	x"078107d1",	x"079207d6",	x"0799075d",	
					x"32607031",	x"07290783",	x"074407a0",	x"072a0771",	
					x"07400780",	x"075f079b",	x"077d079a",	x"075907a2",	
					x"075c077d",	x"077607cc",	x"078e07c3",	x"07b707b5",	
					x"07c307cb",	x"07bf07e2",	x"07dc0814",	x"07d70806",	
					x"07f607d1",	x"07af07ef",	x"07d407fe",	x"07f20809",	
					x"07e1081f",	x"07f70819",	x"07f3081a",	x"07f0082b",	
					x"07fa081b",	x"07e8084c",	x"080b0822",	x"08170823",	
					x"08250862",	x"0821085a",	x"08210870",	x"08350836",	
					x"081f0749",	x"000a0004",	x"f4e55720",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0361002e",	x"07610763",	x"0774074d",	
					x"077a0741",	x"07400748",	x"074c077c",	x"075d0747",	
					x"07570779",	x"075a076d",	x"07a60797",	x"07b20796",	
					x"07a607a0",	x"07b807b7",	x"07ab0795",	x"07b60794",	
					x"07b607bc",	x"0793078b",	x"07a60777",	x"079807a3",	
					x"07b207a4",	x"07a607ab",	x"07a10798",	x"07c20796",	
					x"07bb07b6",	x"0782072c",	x"077d076c",	x"07a507c4",	
					x"079f07a3",	x"07ac07aa",	x"07a307a7",	x"07a4079e",	
					x"07a90792",	x"0765076c",	x"0361102e",	x"076c074d",	
					x"075e0742",	x"07560744",	x"074e0740",	x"073c0742",	
					x"07530778",	x"075a073f",	x"07620750",	x"076f0769",	
					x"07750785",	x"07840794",	x"07940794",	x"07a60780",	
					x"079e0797",	x"079a0789",	x"07590748",	x"076c0756",	
					x"0787076f",	x"07840795",	x"079a0797",	x"07a90787",	
					x"079007a4",	x"07a20768",	x"077e0750",	x"077e078b",	
					x"07940788",	x"07760794",	x"07a507a1",	x"07b00797",	
					x"07900787",	x"079b0799",	x"07870740",	x"0361202e",	
					x"07480746",	x"0747073a",	x"074a071f",	x"072a0724",	
					x"07470730",	x"0751076d",	x"076b0778",	x"07910722",	
					x"07610765",	x"07830760",	x"075b0770",	x"078e078a",	
					x"0773075f",	x"07830757",	x"0772077d",	x"0776072c",	
					x"076a076e",	x"076a0762",	x"07680775",	x"07850772",	
					x"07730777",	x"0780077f",	x"0769075f",	x"0770073d",	
					x"077c0775",	x"0770078c",	x"078b0774",	x"0791078f",	
					x"077e078a",	x"07820786",	x"07640785",	x"0787070c",	
					x"0361302e",	x"070a0715",	x"06ef0717",	x"0721071f",	
					x"07330740",	x"071d0730",	x"0721072e",	x"07390745",	
					x"0755073d",	x"073b0730",	x"074b0743",	x"073e0766",	
					x"07530749",	x"07420773",	x"0778077b",	x"07470754",	
					x"07440728",	x"0745072c",	x"074b074a",	x"0755075b",	
					x"07550774",	x"077f0772",	x"07540766",	x"075a0752",	
					x"0751073f",	x"07640781",	x"0763076b",	x"075f07ae",	
					x"079a07b1",	x"07850789",	x"07770792",	x"07650791",	
					x"07710736",	x"000a0004",	x"4b1a55e8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0362402e",	x"072d073f",	x"07480734",	
					x"07210722",	x"070c0727",	x"0722074f",	x"0755076d",	
					x"07630759",	x"074b072c",	x"07320775",	x"076e0786",	
					x"078e0782",	x"07880787",	x"07820787",	x"07a30785",	
					x"07910780",	x"0781074d",	x"076f079b",	x"07a007b7",	
					x"07a007b5",	x"07ae07c0",	x"07b907bc",	x"07b707a7",	
					x"0798079d",	x"0799077a",	x"079407ac",	x"07b007d0",	
					x"07bf07d4",	x"07d607db",	x"07b907da",	x"07b507d2",	
					x"07a407ce",	x"07aa0797",	x"0362502e",	x"07600784",	
					x"077c07a2",	x"07620765",	x"075f078e",	x"07930780",	
					x"07820785",	x"07870784",	x"07ad078d",	x"078807a7",	
					x"07c207b2",	x"07ab07d8",	x"07e107cc",	x"07ba07e3",	
					x"07e207bb",	x"07a807c5",	x"079e0787",	x"079f07cf",	
					x"07f007bf",	x"079c07d6",	x"07cc07f9",	x"07e307f0",	
					x"07e107e7",	x"07a907db",	x"07d407d2",	x"07b507ef",	
					x"07bd07fe",	x"07bb0808",	x"07ee0813",	x"07ed07ff",	
					x"07ec0808",	x"07d907eb",	x"07da07c1",	x"0362602e",	
					x"078407a2",	x"079e07b7",	x"07820792",	x"078307b9",	
					x"078207c7",	x"07ba07c7",	x"07a907b1",	x"079507ae",	
					x"078e07f6",	x"07d207fc",	x"07cf07ed",	x"07eb07fd",	
					x"07ec07f5",	x"081607eb",	x"07e507e7",	x"07be07c2",	
					x"07c207fa",	x"080207f9",	x"07f00806",	x"07fb0831",	
					x"0802081a",	x"07fa0810",	x"07fd0828",	x"07d10808",	
					x"08070831",	x"0822082f",	x"081b084d",	x"08390846",	
					x"082e084f",	x"082a083d",	x"08220845",	x"080a07be",	
					x"0362702e",	x"079a07c3",	x"07a907d9",	x"07ac07b2",	
					x"079507c8",	x"07cf07cf",	x"07c5082e",	x"080007ff",	
					x"083207f9",	x"07fc082a",	x"08110820",	x"081e0856",	
					x"085f086c",	x"086b0878",	x"085c0860",	x"08550846",	
					x"0849083b",	x"083b0874",	x"0867087c",	x"086d087b",	
					x"085c089e",	x"089008ae",	x"08900896",	x"087e085a",	
					x"08780860",	x"08860886",	x"089108b9",	x"08a208bc",	
					x"08b108bf",	x"08b208aa",	x"08d208d1",	x"08b508bb",	
					x"089306d0",	x"000a0004",	x"7d0691d0",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1363002e",	x"06d806cc",	x"06de06f8",	
					x"070406b9",	x"06ba06e2",	x"06f706ff",	x"07040711",	
					x"070106f0",	x"06fb06e8",	x"06fa06ea",	x"073c072d",	
					x"07270723",	x"07120726",	x"07380722",	x"0727072d",	
					x"0739072c",	x"073f06ee",	x"06fa0709",	x"071f0724",	
					x"071b0719",	x"07300736",	x"0724073e",	x"07300730",	
					x"07180708",	x"071706d6",	x"07200704",	x"071b071d",	
					x"070d0738",	x"0721071b",	x"073a0747",	x"0733074e",	
					x"0741071c",	x"071c06d4",	x"1363102e",	x"06d506d2",	
					x"06dc06cc",	x"06db06c7",	x"06d306c7",	x"06c006fa",	
					x"06f606f6",	x"06f90710",	x"070906d2",	x"07080701",	
					x"07030707",	x"071d0711",	x"07310732",	x"073e06fa",	
					x"0708071c",	x"072a070d",	x"072606c5",	x"06f9070a",	
					x"071d06ff",	x"07100712",	x"072e0719",	x"0718070e",	
					x"071c06fa",	x"0717072c",	x"072806cd",	x"07050727",	
					x"07210729",	x"071b0735",	x"07220723",	x"07370739",	
					x"0763073c",	x"07370727",	x"071a06b8",	x"1363202e",	
					x"06bf06d0",	x"06d406cb",	x"06df06b6",	x"069706b6",	
					x"06cb06c0",	x"06db06d6",	x"06f506dd",	x"06fc06bb",	
					x"06f206f8",	x"0710070a",	x"070f070a",	x"071106fe",	
					x"07070715",	x"070b06f8",	x"06fc0701",	x"070e06c2",	
					x"06d806cf",	x"06da06f6",	x"070c0706",	x"070a0709",	
					x"06f50717",	x"070b071b",	x"06ee070d",	x"070d06e2",	
					x"06fc06e8",	x"06fe0710",	x"0714071b",	x"071e071f",	
					x"071d0720",	x"07280728",	x"07130712",	x"06e806ad",	
					x"1363302e",	x"068506be",	x"069306bf",	x"06ab069e",	
					x"06a406dc",	x"06c206cb",	x"06d906e2",	x"06e906d6",	
					x"06c906c3",	x"06c506c1",	x"06cb06e5",	x"06ef0708",	
					x"06f706fb",	x"06fc06e4",	x"06eb0707",	x"070e06e1",	
					x"06d406c7",	x"06c706d3",	x"06e706f7",	x"06f80702",	
					x"06f7070a",	x"06fb0714",	x"06ff070b",	x"071106ef",	
					x"06f206ec",	x"06f506e7",	x"06ef0701",	x"06f6070e",	
					x"06f60727",	x"06f40723",	x"07080724",	x"07090726",	
					x"06f906d7",	x"000a0004",	x"51c91dae",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"1364402e",	x"06c906d2",	x"06a506e6",	
					x"06d206e6",	x"06d906da",	x"06cd06ea",	x"06e006e8",	
					x"07010701",	x"071d06e0",	x"06d806f9",	x"07100701",	
					x"07160711",	x"07070728",	x"071c0721",	x"07330728",	
					x"071d0728",	x"072c06cb",	x"070e071c",	x"0714070e",	
					x"070f0738",	x"07480746",	x"07410734",	x"072c0737",	
					x"07480737",	x"072a0728",	x"07430740",	x"074d0746",	
					x"074c0756",	x"074c0753",	x"07520763",	x"07610784",	
					x"0752077a",	x"07470703",	x"1364502e",	x"06db0710",	
					x"07080733",	x"070606f7",	x"070d0712",	x"070e0715",	
					x"06fd0750",	x"07380749",	x"07360727",	x"0720074a",	
					x"074b075a",	x"074b074a",	x"075d0763",	x"0755075e",	
					x"0750076a",	x"0751073d",	x"071b072e",	x"0735073c",	
					x"072f0766",	x"07380769",	x"07730783",	x"07500780",	
					x"07610778",	x"075f0785",	x"0745073d",	x"074e0770",	
					x"076507a2",	x"0773078e",	x"07710796",	x"076b07a0",	
					x"0783079b",	x"0782078f",	x"07630716",	x"1364602e",	
					x"06dc071e",	x"071b072e",	x"06fd0719",	x"07160731",	
					x"072b0757",	x"07330754",	x"07400755",	x"072b072d",	
					x"0716076b",	x"077707ad",	x"0784077a",	x"0785078a",	
					x"0781079f",	x"07930784",	x"076d077f",	x"075f0770",	
					x"0752078f",	x"079b0794",	x"078c07ab",	x"07a507d4",	
					x"07ae07c2",	x"079b07ad",	x"079a0799",	x"07960793",	
					x"079707c3",	x"07cd07c2",	x"079b07d8",	x"07c207ef",	
					x"07bc07e5",	x"07c007f2",	x"07ba07cd",	x"07a10736",	
					x"1364702e",	x"07250757",	x"076c0768",	x"07530758",	
					x"07510795",	x"07520781",	x"077e07b8",	x"07c107a7",	
					x"07ae0755",	x"076007ca",	x"07d107e7",	x"07d407f7",	
					x"080e0822",	x"07ed07f1",	x"07f707eb",	x"07ca07ea",	
					x"07de07be",	x"07b107d8",	x"07c307ed",	x"07ce0822",	
					x"08080823",	x"08040836",	x"081d083c",	x"080f080a",	
					x"081f0815",	x"083c0826",	x"0805082c",	x"0819083e",	
					x"0836087a",	x"08310868",	x"083f0875",	x"08520842",	
					x"083d0731",	x"000a0004",	x"86e15cae",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2365002e",	x"073c075a",	x"07550766",	
					x"079c0786",	x"07780788",	x"078c07a5",	x"07bc0798",	
					x"07a6078c",	x"079a0782",	x"078307a4",	x"07b807b0",	
					x"07c707a2",	x"07cf07a1",	x"079f07a7",	x"07a807a2",	
					x"07a90753",	x"078d076b",	x"0783078a",	x"079b078c",	
					x"0797079b",	x"07b6079c",	x"07d0078a",	x"079607cc",	
					x"07dc07b6",	x"0798077f",	x"07ab079e",	x"0786078f",	
					x"07d5079d",	x"079b07cb",	x"07a107d0",	x"07c907bb",	
					x"079507b7",	x"07bd0746",	x"2365102e",	x"074b0752",	
					x"0752073e",	x"07580760",	x"078d0751",	x"07780778",	
					x"0763077a",	x"0788077b",	x"0788074e",	x"0784079b",	
					x"07ae07c1",	x"07b807a0",	x"079f0769",	x"07980767",	
					x"07970787",	x"07a70756",	x"07a10754",	x"07750776",	
					x"07940777",	x"07890791",	x"07920777",	x"07870778",	
					x"079f0795",	x"078e07a6",	x"07bb0749",	x"07a0078b",	
					x"0794079b",	x"07ab07ac",	x"07a10779",	x"07bb07ac",	
					x"07ad07bc",	x"07b507a3",	x"079b0741",	x"2365202e",	
					x"07430748",	x"07280720",	x"073a0713",	x"0741071b",	
					x"07610754",	x"07830765",	x"0786075b",	x"07790759",	
					x"0763075c",	x"077a0761",	x"076a0772",	x"07750770",	
					x"07810777",	x"078f0775",	x"078a0770",	x"076a072e",	
					x"072e0779",	x"07750777",	x"07690776",	x"0780075d",	
					x"07680764",	x"077e0770",	x"076e074e",	x"0756073a",	
					x"076a0784",	x"07690774",	x"07690771",	x"0770076b",	
					x"07720780",	x"078b078c",	x"077d079e",	x"078906ea",	
					x"2365302e",	x"06fb0708",	x"0709073a",	x"070a073b",	
					x"073b0735",	x"0757072d",	x"073b0735",	x"072b0731",	
					x"072c071e",	x"073a075e",	x"0745076c",	x"076c075b",	
					x"07670773",	x"07590763",	x"077b074c",	x"075d076a",	
					x"07510716",	x"07280736",	x"07530756",	x"07580772",	
					x"074b0774",	x"0753076b",	x"07640771",	x"07530765",	
					x"07500750",	x"074e077a",	x"07510775",	x"07690775",	
					x"07680798",	x"0771079a",	x"076c0783",	x"0764079c",	
					x"076c0718",	x"000a0004",	x"cee1586e",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"2366402e",	x"070a0729",	x"07240751",	
					x"07360745",	x"073c073e",	x"075b073e",	x"07590752",	
					x"07350737",	x"07540744",	x"07590759",	x"07760774",	
					x"0781077c",	x"07a0077f",	x"0780076f",	x"07790775",	
					x"07890770",	x"077c076e",	x"077b076b",	x"07820773",	
					x"07960768",	x"07b507b9",	x"07a407b2",	x"07b1079a",	
					x"07b2079d",	x"07b20796",	x"07b60797",	x"07a60796",	
					x"07a2079c",	x"07a307b5",	x"07ca07c1",	x"07d307bb",	
					x"07c407b7",	x"07c60735",	x"2366502e",	x"0726075f",	
					x"07700768",	x"07700768",	x"07720798",	x"077e078f",	
					x"079c07b2",	x"07af07a2",	x"07b907b1",	x"07b307cd",	
					x"07c507d1",	x"07ce07c8",	x"07d207b6",	x"07bf07cc",	
					x"07b407c1",	x"07b307ba",	x"07bd0796",	x"079207c3",	
					x"07ba07c6",	x"07a207d1",	x"07b70813",	x"07ba0805",	
					x"07d107d5",	x"07d007e3",	x"07da07d3",	x"07df07d5",	
					x"07a907f2",	x"07dc07fa",	x"07e70808",	x"07d60814",	
					x"07ee080c",	x"07e30808",	x"07da074c",	x"2366602e",	
					x"073a076e",	x"075e07b9",	x"0781077b",	x"07810791",	
					x"079007a4",	x"079d07ad",	x"07bc078d",	x"07a407c7",	
					x"07d907fe",	x"07f607f3",	x"07e307f3",	x"07f40804",	
					x"07e40807",	x"07f80806",	x"07e907e8",	x"07c807d3",	
					x"07b007d6",	x"07e907fb",	x"07e2080b",	x"07fc0815",	
					x"07ee0818",	x"080c0809",	x"08090815",	x"08040802",	
					x"0810082f",	x"08170823",	x"08100840",	x"08240864",	
					x"0822085b",	x"08220853",	x"08220834",	x"081507c4",	
					x"2366702e",	x"077107ba",	x"07ad07da",	x"07b507cc",	
					x"07c607f2",	x"07d30816",	x"0816083c",	x"082f07ce",	
					x"07ee07fb",	x"081f0877",	x"0849085c",	x"0852083a",	
					x"08220850",	x"08390852",	x"08480868",	x"08320831",	
					x"0831083f",	x"0834085c",	x"08580879",	x"085f0868",	
					x"085c0884",	x"08610871",	x"08920886",	x"087f087a",	
					x"085b0869",	x"08940888",	x"089208a6",	x"087c08a7",	
					x"088608f9",	x"087a08da",	x"08a508db",	x"08c908bd",	
					x"089806e7",	x"000a0004",	x"fc808f1b",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3367002e",	x"06e3069e",	x"06a806ab",	
					x"06c906b2",	x"06ab06fe",	x"06f406d1",	x"06ff06f3",	
					x"070a06d9",	x"06f606eb",	x"06e106e0",	x"071f06f8",	
					x"071d0702",	x"074f0729",	x"072606f6",	x"071006f4",	
					x"070a06c7",	x"06d606e4",	x"06ec06ff",	x"070a06fc",	
					x"071206fc",	x"070306ff",	x"07090707",	x"070f06ff",	
					x"06f5071a",	x"072106f9",	x"071b06d5",	x"06f90724",	
					x"071906f6",	x"070f06eb",	x"06fc06f6",	x"071f0720",	
					x"06fb071e",	x"06ff06c8",	x"3367102e",	x"06bb06b7",	
					x"06d406ab",	x"06c40695",	x"06c606cb",	x"06d006e1",	
					x"06db06e0",	x"06da06e4",	x"06ec06d6",	x"06f0070a",	
					x"06fe0731",	x"07260707",	x"070106f3",	x"070806d9",	
					x"06e406d2",	x"06eb06ba",	x"06ba06d1",	x"06e106e1",	
					x"070406dc",	x"070806f5",	x"070b06f4",	x"070e06f8",	
					x"07200718",	x"071e06ea",	x"06f906d3",	x"06e30703",	
					x"070806fa",	x"06f7070a",	x"071006eb",	x"06f30706",	
					x"0707072a",	x"0719071f",	x"0718069d",	x"3367202e",	
					x"06940687",	x"06a006a6",	x"06b806bf",	x"06c306b4",	
					x"06bb06c2",	x"06da06bb",	x"06d206a9",	x"06db06c5",	
					x"06e406f4",	x"070e06ef",	x"070106f1",	x"06f206e2",	
					x"06f006dd",	x"06e406d8",	x"06bf06c7",	x"06d106ab",	
					x"06b406e8",	x"06dd06cf",	x"06df06d8",	x"06e606d0",	
					x"06de06c4",	x"06c706d5",	x"06d106e5",	x"06ed06dc",	
					x"06fd06e2",	x"06f206fb",	x"06f906d6",	x"06df06f8",	
					x"070506dd",	x"06dd06fa",	x"06e10708",	x"06e906a3",	
					x"3367302e",	x"068f06ac",	x"06aa0696",	x"06a5066a",	
					x"068b06b2",	x"069006a3",	x"06d206da",	x"06c206a0",	
					x"069d068c",	x"06a206d4",	x"06cd06c2",	x"06c006d4",	
					x"06cd06cb",	x"06d006c4",	x"06b706c5",	x"06b206db",	
					x"06c306a1",	x"06a706dd",	x"06dc06d6",	x"06e206e8",	
					x"071306f0",	x"06d806de",	x"06f106fc",	x"06dc06da",	
					x"06cd06d5",	x"06ce06f8",	x"06e906e5",	x"06b006ff",	
					x"06eb06f8",	x"06df0706",	x"06e8070b",	x"06e6070b",	
					x"06e306a5",	x"000a0004",	x"c4670ec3",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3368402e",	x"068806ae",	x"069d06b1",	
					x"06a906cf",	x"06c606cd",	x"06bc06ac",	x"06ac06c4",	
					x"06b406d4",	x"06d806cf",	x"06d706dd",	x"070306fc",	
					x"06fa06f6",	x"070006f8",	x"06f106f7",	x"070a06e0",	
					x"06fd06e4",	x"06f106d4",	x"06f806f1",	x"06f106f9",	
					x"07190707",	x"07160703",	x"07150715",	x"0718070d",	
					x"07140731",	x"0727070e",	x"070d0712",	x"0726070c",	
					x"0710072c",	x"072f073a",	x"072f073a",	x"072f073a",	
					x"073c074b",	x"072d06cc",	x"3368502e",	x"06d806cf",	
					x"06be06e0",	x"06ad06e7",	x"06d206ea",	x"06e106f3",	
					x"06cd0709",	x"06fc0719",	x"071806fb",	x"06f2072f",	
					x"072b0727",	x"07430729",	x"0743071b",	x"0726071d",	
					x"0722071c",	x"07180709",	x"071106fb",	x"070d0723",	
					x"071f0731",	x"071d072c",	x"07200738",	x"07290749",	
					x"07160749",	x"0727073f",	x"0713074a",	x"072b075f",	
					x"072d0752",	x"072f0766",	x"07370765",	x"0740075d",	
					x"07450771",	x"07400769",	x"074a06c4",	x"3368602e",	
					x"06bd06e0",	x"06be06f1",	x"06e006fa",	x"06ed0703",	
					x"06f006ec",	x"06e7073c",	x"07260715",	x"07070721",	
					x"07020741",	x"0742075f",	x"072e074a",	x"072f0759",	
					x"0757074c",	x"07370754",	x"07450746",	x"074f071f",	
					x"0720076a",	x"07560748",	x"074f0761",	x"074e0780",	
					x"07600774",	x"07840777",	x"0766077d",	x"0767076c",	
					x"077e0770",	x"0776079e",	x"0778078c",	x"076807a6",	
					x"077907a8",	x"077f07aa",	x"078907b9",	x"076a0717",	
					x"3368702e",	x"071d074d",	x"072d0724",	x"0738072a",	
					x"0721074e",	x"072b071c",	x"07310760",	x"07540763",	
					x"0750077a",	x"077b07aa",	x"079e07cf",	x"07a50790",	
					x"077e07ce",	x"07b107c2",	x"07ac07f3",	x"07880791",	
					x"07a3079a",	x"07b307c4",	x"079c07d6",	x"07ac07cb",	
					x"07c407f4",	x"07dc07d2",	x"07dc07ee",	x"07dc07f1",	
					x"07cc07a5",	x"07ab07de",	x"07e307de",	x"07e80830",	
					x"07f00836",	x"07da0830",	x"081e082c",	x"0822081b",	
					x"0813079c",	x"000a0004",	x"eed34427",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"0369002f",	x"078a0790",	x"07a70792",	
					x"077e0792",	x"078407bc",	x"07930762",	x"07620762",	
					x"076e076f",	x"078b0766",	x"0791078f",	x"07a107a2",	
					x"07ba07c0",	x"07c607af",	x"07c907b0",	x"07da07d2",	
					x"07c207bf",	x"07ca078b",	x"078d078f",	x"07a2079c",	
					x"07b807a5",	x"079e07a5",	x"07b0079a",	x"07a2079b",	
					x"07a9078a",	x"07af077f",	x"07ae07c8",	x"07bf07b2",	
					x"079a07ba",	x"07bf07b1",	x"07b307c4",	x"07bb07bf",	
					x"07b107c3",	x"07a10771",	x"0369102f",	x"0794077d",	
					x"07720775",	x"079f0769",	x"075a074c",	x"0741074e",	
					x"07490724",	x"07490735",	x"075c075e",	x"077c078e",	
					x"0797079c",	x"07ab07bc",	x"07ac0798",	x"07a50790",	
					x"07b70787",	x"078a0783",	x"078b0775",	x"078b078f",	
					x"07aa07b4",	x"07bf079f",	x"078e07bc",	x"07a40781",	
					x"078d079f",	x"078107ad",	x"079c076e",	x"079d079d",	
					x"07c907a4",	x"07ae07b6",	x"07cb079f",	x"07a707de",	
					x"07ca07d0",	x"07bd07b9",	x"079c0784",	x"0369202f",	
					x"075f0764",	x"0777075d",	x"077f0757",	x"0755073a",	
					x"0752075d",	x"07500749",	x"07420758",	x"07760756",	
					x"075e077c",	x"079c0775",	x"077b077a",	x"07a60777",	
					x"078e0789",	x"0779075e",	x"0761076c",	x"07640737",	
					x"076c0759",	x"07650781",	x"07800792",	x"079c078b",	
					x"077f076c",	x"07780792",	x"078c07a2",	x"07950779",	
					x"0785078a",	x"07830785",	x"077d078b",	x"07a707ac",	
					x"0798079d",	x"079c079a",	x"07760797",	x"07ab0758",	
					x"0369302f",	x"0756074e",	x"0745074d",	x"07550763",	
					x"0756076b",	x"07430754",	x"07320761",	x"074e0750",	
					x"074d0745",	x"0732077c",	x"0765078b",	x"074f0794",	
					x"0776078e",	x"07820797",	x"07960787",	x"07810786",	
					x"07720746",	x"0751079e",	x"078a0792",	x"077707a2",	
					x"0785078e",	x"076707a2",	x"079007b9",	x"079807b1",	
					x"0783078b",	x"077707b3",	x"0784079c",	x"076407c4",	
					x"07a607ca",	x"07a307b5",	x"079907cf",	x"07a407dc",	
					x"07a70794",	x"000a0004",	x"566f650b",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"036a402f",	x"076d078f",	x"0787076a",	
					x"07650774",	x"07460780",	x"07430765",	x"0779079e",	
					x"07a20783",	x"075d078e",	x"07570786",	x"076f07b3",	
					x"079207c5",	x"07af07c8",	x"07a807c7",	x"07ba07c2",	
					x"07ae07bb",	x"07a207b6",	x"07c907c8",	x"07c707e9",	
					x"07cf07ce",	x"07ce07fc",	x"07d607fb",	x"07d207f7",	
					x"07c40801",	x"07d50804",	x"07c50804",	x"07e50825",	
					x"07f0082b",	x"08020821",	x"07ef0814",	x"07fa0844",	
					x"07f8084d",	x"080d07f6",	x"036a502f",	x"0790079f",	
					x"07a307a7",	x"079b07c8",	x"07bf07c6",	x"078807c8",	
					x"07c507c6",	x"078107ea",	x"07d507ff",	x"07cc07f3",	
					x"07f407e5",	x"07fa0809",	x"080807ff",	x"07d20802",	
					x"07f1080c",	x"07f1080f",	x"07f107eb",	x"07bc0809",	
					x"07db07f0",	x"07b60804",	x"07d40810",	x"07d60817",	
					x"07f6083f",	x"07f3082f",	x"07f70806",	x"07e7087d",	
					x"08150853",	x"080e0860",	x"081d0887",	x"08110868",	
					x"082a0861",	x"08110858",	x"082207fe",	x"036a602f",	
					x"07cc07df",	x"07b20815",	x"07bf07d9",	x"07ae07fc",	
					x"07b407e4",	x"07bf07c7",	x"07b0081d",	x"07ce0829",	
					x"07dd0812",	x"07ed083a",	x"07ef0821",	x"07d20818",	
					x"07fc0820",	x"07f60833",	x"07f2083a",	x"07f60844",	
					x"07f30838",	x"080c0855",	x"08190832",	x"082b085e",	
					x"08140867",	x"0817085d",	x"0813086d",	x"081e0864",	
					x"082d0871",	x"0822088b",	x"083e089d",	x"086408b6",	
					x"084d08bb",	x"085308b3",	x"087008af",	x"088107f0",	
					x"036a702f",	x"07b50828",	x"07de0800",	x"07af0803",	
					x"07b9081e",	x"077c07e9",	x"0790081d",	x"07b80815",	
					x"07fb0800",	x"07fb0857",	x"0820084a",	x"08300886",	
					x"0867088b",	x"086408ad",	x"087208aa",	x"08570892",	
					x"08640876",	x"083908ba",	x"086608cc",	x"085d08c3",	
					x"087808d1",	x"088508ed",	x"08ce08e2",	x"086f08bb",	
					x"088f08ca",	x"08a708c8",	x"088f0909",	x"08a30905",	
					x"090108fd",	x"08bc08f6",	x"08c30927",	x"08db090d",	
					x"08e806f9",	x"000a0004",	x"8de6b473",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"136b002f",	x"070d0711",	x"07210717",	
					x"071206f0",	x"06fa0709",	x"06e306ec",	x"06f806f1",	
					x"06e006bd",	x"06d906d3",	x"06d506db",	x"06f8071c",	
					x"07200724",	x"073606f8",	x"07220734",	x"07430755",	
					x"075b06ff",	x"071b06ed",	x"071b0718",	x"072e072f",	
					x"07270719",	x"073a0723",	x"0733072e",	x"074b0729",	
					x"072e071b",	x"073006f3",	x"07030721",	x"0741073d",	
					x"07390740",	x"072c0710",	x"07200740",	x"07270745",	
					x"0738071d",	x"07150705",	x"136b102f",	x"06c806c9",	
					x"06e006ca",	x"06ee06c5",	x"06dd06d0",	x"06ca06d1",	
					x"06c206c5",	x"06d106d6",	x"06af06a6",	x"06b90708",	
					x"071a070e",	x"070506ec",	x"072c0728",	x"073b0716",	
					x"07290713",	x"072b0709",	x"071806ed",	x"06fd0706",	
					x"0707071e",	x"0732071c",	x"071a071c",	x"071e0718",	
					x"071d072b",	x"072b0724",	x"071106e8",	x"07080724",	
					x"07130734",	x"07270744",	x"0750072b",	x"073c073c",	
					x"072e0759",	x"07470738",	x"073406e3",	x"136b202f",	
					x"06e706fb",	x"06fb06e2",	x"06f106f3",	x"070606de",	
					x"06a106d5",	x"06f606df",	x"070a06af",	x"06ee06ba",	
					x"06ef06c0",	x"06fa06f0",	x"07190719",	x"07130714",	
					x"071d06f5",	x"06f406f1",	x"07030723",	x"070b06e0",	
					x"06f106ee",	x"070306dd",	x"06fd0709",	x"070f071d",	
					x"06f90713",	x"070b0709",	x"07010717",	x"070606d5",	
					x"071f06f9",	x"07140723",	x"071b0712",	x"07150714",	
					x"06f30720",	x"072d071d",	x"07060720",	x"06f706d2",	
					x"136b302f",	x"06bf06d5",	x"06be06e3",	x"06cc06c0",	
					x"06c006bb",	x"06a906e9",	x"06ae06b8",	x"06b806aa",	
					x"06b006a1",	x"06ac06de",	x"06d306ef",	x"06e4071d",	
					x"07000719",	x"06d1070d",	x"0713070d",	x"06ed06f5",	
					x"06df06ee",	x"06e60709",	x"06fe070a",	x"070d070f",	
					x"070d0733",	x"071e072d",	x"07020718",	x"07000726",	
					x"071c06f2",	x"06f9070e",	x"06f40747",	x"070d0746",	
					x"07140747",	x"071a0743",	x"071e073a",	x"07170739",	
					x"071a06e4",	x"000a0004",	x"544521d8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"136c402f",	x"06ad06c9",	x"06c906f4",	
					x"06d006fc",	x"06f80702",	x"06d606f9",	x"06db06d4",	
					x"06d106e1",	x"06f106ef",	x"06e20749",	x"07150739",	
					x"0725072f",	x"07270731",	x"07200739",	x"073f0743",	
					x"071e074a",	x"0748072d",	x"0718073b",	x"07420752",	
					x"074e0756",	x"074d0767",	x"0751073c",	x"07420759",	
					x"07480743",	x"0735074c",	x"074e0796",	x"076e076e",	
					x"07540761",	x"075b0773",	x"07650784",	x"07750792",	
					x"07680782",	x"0730073b",	x"136c502f",	x"06ff0731",	
					x"07150715",	x"06da071a",	x"07000712",	x"06f00730",	
					x"06fd0752",	x"06e20744",	x"07180707",	x"07130782",	
					x"074f0761",	x"073a0779",	x"07560775",	x"07680767",	
					x"075c0775",	x"0756076a",	x"07460749",	x"073e0787",	
					x"07650795",	x"07710792",	x"077a07ac",	x"076807a6",	
					x"077b0795",	x"075b078d",	x"075d0796",	x"078e07b3",	
					x"079307d0",	x"078507b9",	x"079307ad",	x"078b07d8",	
					x"079407cb",	x"078e079b",	x"0764073a",	x"136c602f",	
					x"06f8074a",	x"0724074d",	x"07320739",	x"071b074e",	
					x"071d0769",	x"06f80757",	x"074e075b",	x"0727074d",	
					x"0712076e",	x"077d0777",	x"07720780",	x"078007ad",	
					x"077f07b4",	x"078807b2",	x"078607a6",	x"079307a2",	
					x"078507b8",	x"079e07ca",	x"07a907fd",	x"07b107cb",	
					x"07a707d3",	x"079907d8",	x"079d07cd",	x"07af07c0",	
					x"07a307e1",	x"07b707f0",	x"07a507f3",	x"07b007fe",	
					x"07c407ec",	x"07d307f4",	x"07bd07d7",	x"07b2075c",	
					x"136c702f",	x"07120779",	x"076f07bc",	x"076b0775",	
					x"075007a4",	x"07260797",	x"074c0783",	x"07410781",	
					x"075507bd",	x"077907b7",	x"079a07e0",	x"07b207f8",	
					x"07ec082a",	x"07ee081d",	x"08010830",	x"07ec082c",	
					x"07bf07ff",	x"07bd0827",	x"080d086b",	x"081a083f",	
					x"08110832",	x"08160846",	x"080e0856",	x"0821081c",	
					x"084d080d",	x"0823084f",	x"084b0881",	x"080a0879",	
					x"08410870",	x"0830088d",	x"085108a9",	x"08450856",	
					x"081c0763",	x"000a0004",	x"89d86b7a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"236d002f",	x"075a0774",	x"075d078d",	
					x"078f0761",	x"0770078b",	x"0764075e",	x"075a0787",	
					x"076c0776",	x"07840782",	x"078a07b9",	x"07b707c6",	
					x"07c807cb",	x"07c107b0",	x"07af07a4",	x"07a4079b",	
					x"079407a3",	x"07a00769",	x"078307ac",	x"07ca07a7",	
					x"07b507be",	x"07bd079c",	x"07a507a9",	x"0798078b",	
					x"07ad07bb",	x"079d07bb",	x"07cc0798",	x"07b607b7",	
					x"07bc07d7",	x"07be07cd",	x"079707a3",	x"07b307dd",	
					x"079a0796",	x"07890765",	x"236d102f",	x"07680757",	
					x"07550752",	x"076b0740",	x"073f0720",	x"0749076f",	
					x"0768075c",	x"076f0755",	x"0769075b",	x"0744079d",	
					x"079e07a4",	x"0799078f",	x"079e0781",	x"078e0784",	
					x"07900788",	x"07af078a",	x"07bf0747",	x"075c076a",	
					x"07aa07a5",	x"07b1078b",	x"07a90799",	x"07b60794",	
					x"07b507a6",	x"07ac0792",	x"079b0757",	x"07b9078d",	
					x"07ae07a5",	x"07bc07b2",	x"07a307a1",	x"07ab07ab",	
					x"079e07c9",	x"079d07a0",	x"07bc0708",	x"236d202f",	
					x"071f0727",	x"07300746",	x"076c0753",	x"07630745",	
					x"073b0732",	x"07410762",	x"07790768",	x"07660726",	
					x"073a076b",	x"078e0780",	x"077a0770",	x"07870767",	
					x"078d0784",	x"0784078b",	x"078307a5",	x"0773076f",	
					x"076e0782",	x"07860787",	x"07520785",	x"07860768",	
					x"0778078d",	x"07900789",	x"07980797",	x"07860787",	
					x"07840787",	x"0782077d",	x"07870790",	x"079c0773",	
					x"0786078c",	x"078207d3",	x"07900793",	x"07710737",	
					x"236d302f",	x"071d0723",	x"07250732",	x"0728072c",	
					x"073d072f",	x"07130721",	x"072e074a",	x"07280755",	
					x"07340718",	x"07470747",	x"07580753",	x"075d0769",	
					x"076c0769",	x"0751073f",	x"0747074c",	x"07660751",	
					x"075a073e",	x"0745076f",	x"07630766",	x"07660778",	
					x"075f076e",	x"075e0779",	x"0767079b",	x"07610777",	
					x"07600771",	x"076407ce",	x"07670795",	x"0770078d",	
					x"07690794",	x"075f07a4",	x"077c0799",	x"077e0796",	
					x"07690734",	x"000a0004",	x"cfe05dcb",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"236e402f",	x"07220757",	x"07410731",	
					x"071a0747",	x"073b075c",	x"073e075c",	x"07560763",	
					x"07470763",	x"0757076d",	x"074f0785",	x"078d0785",	
					x"078b078f",	x"0790079a",	x"078a0796",	x"0794078d",	
					x"0797079b",	x"078c079f",	x"079d07c5",	x"07c307b3",	
					x"07b007cf",	x"079b07ca",	x"07a207c3",	x"07d007bd",	
					x"07cf07b5",	x"07c507b7",	x"07c907d1",	x"07bf07cf",	
					x"07c907d4",	x"07e007c0",	x"07d007e9",	x"07d807df",	
					x"07cb07c9",	x"07c00769",	x"236e502f",	x"073b076a",	
					x"07620777",	x"0737079b",	x"077f07a8",	x"077607a8",	
					x"0783077d",	x"077407d6",	x"07c307ac",	x"079407b9",	
					x"07b407e1",	x"07c807d0",	x"07c007e2",	x"07b60805",	
					x"07c907dd",	x"07c707da",	x"07b807e3",	x"07b907ff",	
					x"07d80801",	x"07b807f6",	x"07d9081b",	x"07e90821",	
					x"07fb080f",	x"07f10842",	x"08070803",	x"07fe081f",	
					x"07dc0818",	x"07dd0826",	x"07de083d",	x"07d70849",	
					x"07fb083d",	x"07ff0821",	x"07e8077f",	x"236e602f",	
					x"07720784",	x"076907c8",	x"07800799",	x"078a07ab",	
					x"075c07cb",	x"076607da",	x"07b607e5",	x"07c40802",	
					x"07bd082b",	x"07cc0829",	x"07e80829",	x"08030852",	
					x"07eb081b",	x"07f60825",	x"07f10829",	x"07d90809",	
					x"07ea0847",	x"080e0828",	x"07e90833",	x"07fe0853",	
					x"0812085a",	x"08130846",	x"08180866",	x"080c0849",	
					x"082a083d",	x"081e0837",	x"08180867",	x"082f0873",	
					x"08310873",	x"0829087c",	x"083d0862",	x"081307e6",	
					x"236e702f",	x"078007e0",	x"079d07da",	x"078907e8",	
					x"07a107fe",	x"07c607f8",	x"07ea082c",	x"07d30842",	
					x"07f707f3",	x"07d0084c",	x"0817086d",	x"082d088b",	
					x"084f0895",	x"082c08b6",	x"086308a1",	x"085f0878",	
					x"083c087d",	x"083d087c",	x"084f088d",	x"085a0881",	
					x"088508c3",	x"089908ba",	x"088b08cf",	x"089708c3",	
					x"08ab0894",	x"088e08a9",	x"08b608bb",	x"08b308b1",	
					x"08b708ec",	x"089008f0",	x"08bf08f6",	x"08ae08d6",	
					x"08d30703",	x"000a0004",	x"00baa23a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"336f002f",	x"06ec06da",	x"06f806dd",	
					x"06ce06cf",	x"06dc06c9",	x"06cb06f3",	x"06fc06ff",	
					x"06d706af",	x"06ca06f2",	x"06d5070d",	x"072706f8",	
					x"071f06fc",	x"07270720",	x"07390707",	x"073c071a",	
					x"073006fb",	x"06f406d7",	x"06fc071c",	x"06f206e6",	
					x"070506fd",	x"07090701",	x"070b0707",	x"071e071c",	
					x"0727070f",	x"072106d9",	x"070d0708",	x"071c0723",	
					x"072306f9",	x"06f906e6",	x"070606e7",	x"07170704",	
					x"070006f7",	x"06f906bc",	x"336f102f",	x"06c906cc",	
					x"06bf06bd",	x"06c306bb",	x"06ce06bb",	x"06bd06b8",	
					x"06b406c2",	x"06c606c8",	x"06c5069a",	x"06c90702",	
					x"06fe0728",	x"070706fd",	x"070406ee",	x"070206fb",	
					x"06e00700",	x"06f806ff",	x"06f206e1",	x"06c906fa",	
					x"070a06ef",	x"070e06ee",	x"06e406eb",	x"06f806d3",	
					x"06f7070b",	x"07110714",	x"070506ef",	x"06fb0725",	
					x"07250700",	x"071306fe",	x"071806e7",	x"06fd0708",	
					x"0719071a",	x"070a0720",	x"072506c2",	x"336f202f",	
					x"06b306b6",	x"06b606ae",	x"068a06c6",	x"06b00690",	
					x"06990681",	x"06a90690",	x"06a30681",	x"06b706b1",	
					x"06cc06e1",	x"06f306e9",	x"06f706e7",	x"06e606f1",	
					x"06ec06d6",	x"06fe06de",	x"06bf06e9",	x"06df06bf",	
					x"06d10702",	x"06f906e3",	x"06e006eb",	x"06f306e7",	
					x"06e306dd",	x"06e406e8",	x"06f706e3",	x"06ea06cc",	
					x"06f006e6",	x"06ee06e2",	x"06ef06fb",	x"06f306f1",	
					x"06e306e3",	x"06f40707",	x"06f10704",	x"06ea06ca",	
					x"336f302f",	x"069b06b1",	x"069d06b0",	x"06880680",	
					x"068506a6",	x"06830697",	x"068e0695",	x"06a406b2",	
					x"06a906ab",	x"06bb06d4",	x"06c406e0",	x"06c306da",	
					x"06d106df",	x"06d306e8",	x"06c806e6",	x"06c206e1",	
					x"06d306d0",	x"06b206ce",	x"06e406d7",	x"06e206f1",	
					x"0708070e",	x"06fb06e3",	x"06f20709",	x"06d8070e",	
					x"06ce06f3",	x"06d40708",	x"0710070f",	x"06f10714",	
					x"06d80704",	x"06d80710",	x"06de0703",	x"06de06f3",	
					x"06d706b1",	x"000a0004",	x"c47c11c2",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"3370402f",	x"068406b8",	x"06a106b3",	
					x"068006ce",	x"06af06d1",	x"06ac06cb",	x"06a706d3",	
					x"06ae06e8",	x"06b906ed",	x"06ef06f9",	x"06ee070e",	
					x"06ec06ef",	x"06ee06e6",	x"06e10704",	x"06ed0709",	
					x"07150723",	x"071106e5",	x"070d0725",	x"0708072a",	
					x"07360727",	x"07280721",	x"070d0731",	x"0725072c",	
					x"07280743",	x"07370740",	x"072d075f",	x"07380742",	
					x"07370744",	x"07360749",	x"073b0785",	x"07400742",	
					x"07380749",	x"072a0702",	x"3370502f",	x"06df0705",	
					x"06fb0703",	x"06ba06e2",	x"06e6071d",	x"07030710",	
					x"06df072d",	x"07060720",	x"06f40712",	x"070f0731",	
					x"07280740",	x"0739074f",	x"0758074f",	x"073e0758",	
					x"07380754",	x"071c073f",	x"073f0723",	x"07140745",	
					x"07320756",	x"073a0758",	x"073f0772",	x"073c077c",	
					x"072f0785",	x"07520789",	x"0753075c",	x"074107ab",	
					x"075b075d",	x"07380781",	x"074a0787",	x"073e0793",	
					x"076407ab",	x"0763077a",	x"074f0712",	x"3370602f",	
					x"06f70729",	x"06f10721",	x"06d506e5",	x"06db073a",	
					x"06ec071b",	x"07000732",	x"071e0736",	x"07270739",	
					x"071b0761",	x"0746077a",	x"075a077c",	x"074e078e",	
					x"0772077c",	x"07610780",	x"07720778",	x"074b0770",	
					x"07380791",	x"0789079a",	x"07790784",	x"07780798",	
					x"07860789",	x"077e07a6",	x"076f07a4",	x"07a207a4",	
					x"077b07bb",	x"07a007bb",	x"077807c5",	x"077c07b9",	
					x"077b07c5",	x"078d07ac",	x"079507b4",	x"077a072b",	
					x"3370702f",	x"07010746",	x"07070743",	x"07020742",	
					x"07000751",	x"0718075c",	x"0727075f",	x"074207a1",	
					x"075e0775",	x"076907aa",	x"079b07d4",	x"078107ca",	
					x"078f07df",	x"078807e5",	x"07ab07ce",	x"07a107db",	
					x"07bd07ab",	x"077707f7",	x"07c90814",	x"07b307c4",	
					x"07bb07d0",	x"07c407d7",	x"07ca0823",	x"07de0833",	
					x"07dd07ef",	x"07e7083a",	x"07f5083c",	x"07d90835",	
					x"07d20820",	x"07ea0854",	x"07fa0854",	x"08170823",	
					x"07ff0787",	x"000a0004",	x"f3a1548a",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"03710030",	x"07d10799",	x"07ba0785",	
					x"07930786",	x"076e07a8",	x"07b207a9",	x"07ee07e2",	
					x"07f807d7",	x"07e607b5",	x"07d607be",	x"07a807bd",	
					x"081207bf",	x"07d907bf",	x"07d907b4",	x"07f907ca",	
					x"07dd07cd",	x"07e7077c",	x"07b2078d",	x"07de07a9",	
					x"07db07ab",	x"07d007da",	x"07d907d8",	x"081907d1",	
					x"07e407bc",	x"07d60770",	x"079107bb",	x"07c307ff",	
					x"07c507d3",	x"07fe0804",	x"07e10802",	x"07f507ea",	
					x"07d807ee",	x"07f207a2",	x"03711030",	x"080f07a8",	
					x"07c407a3",	x"07be07a9",	x"07bc07bb",	x"07aa07e8",	
					x"07f807df",	x"07e507f0",	x"080807d2",	x"07ff07da",	
					x"07ca07da",	x"07e907d9",	x"080a07fe",	x"080d07ea",	
					x"07e707d9",	x"07d507d7",	x"07e207c8",	x"07b107b6",	
					x"07fc07d7",	x"081307fc",	x"07f907f2",	x"080007fa",	
					x"080607e9",	x"07dc0805",	x"07f40760",	x"07b807c6",	
					x"07d207eb",	x"07f107f8",	x"07ff07f7",	x"07f50811",	
					x"07fc080d",	x"080807ec",	x"07c707a1",	x"03712030",	
					x"07dc0799",	x"079a077d",	x"07a8078e",	x"07c70782",	
					x"07ec07db",	x"07ea07dc",	x"07e607d8",	x"07d907a3",	
					x"07cd07bd",	x"07d007ae",	x"07c507b1",	x"07de07ca",	
					x"07d807bc",	x"07dd07ce",	x"07d507c1",	x"079f075b",	
					x"079d07a8",	x"07e407b6",	x"079a07be",	x"07cf07c1",	
					x"07bb07bf",	x"07d007c3",	x"07bc07c6",	x"07c70771",	
					x"07a107d3",	x"07d407d9",	x"07d807ca",	x"07e707e1",	
					x"07e307e0",	x"07e307c4",	x"079f07e1",	x"07e40734",	
					x"03713030",	x"07720736",	x"07290735",	x"073c0757",	
					x"0762075b",	x"07390756",	x"078d0780",	x"07950782",	
					x"079b0771",	x"07760793",	x"079e079c",	x"07890795",	
					x"07870785",	x"078c0791",	x"0787078f",	x"07680777",	
					x"076c0742",	x"07720782",	x"07a6078d",	x"07a70794",	
					x"078d07a8",	x"07ab07bd",	x"07a307bd",	x"07ab079a",	
					x"075e0732",	x"077b07ae",	x"079407af",	x"07a407da",	
					x"07c407d6",	x"07a207b6",	x"079207d8",	x"07ae07e0",	
					x"07a30781",	x"000a0004",	x"73977aae",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"03724030",	x"0796076c",	x"075e074f",	
					x"0736075c",	x"076b0790",	x"078d0780",	x"07a907a3",	
					x"07aa0798",	x"07940794",	x"078807b7",	x"07aa07b6",	
					x"07cb07be",	x"07c607b8",	x"07bc07b7",	x"07c807b7",	
					x"07ca07ac",	x"07bf079d",	x"079d07ac",	x"07c407ab",	
					x"07ae07db",	x"07df07f7",	x"07f30800",	x"07e007dd",	
					x"07cf0791",	x"07960799",	x"07a807cb",	x"07d9080e",	
					x"07e1080f",	x"08120821",	x"07df0800",	x"07fa0807",	
					x"07e4082d",	x"07ec07da",	x"03725030",	x"07bf07a0",	
					x"07a7079b",	x"077c07b7",	x"07a607cc",	x"07c107c1",	
					x"07e207ef",	x"07e807cf",	x"07e107cd",	x"07de07e4",	
					x"07ff07ed",	x"07e307ff",	x"07f607fe",	x"080d0826",	
					x"082b07cb",	x"07c907d8",	x"07cf07db",	x"07d907e3",	
					x"07dd0808",	x"07de0818",	x"0810081c",	x"08010827",	
					x"080c0830",	x"07f7081a",	x"07e00805",	x"07e90821",	
					x"07f50822",	x"08020842",	x"081d087a",	x"08290849",	
					x"08200852",	x"0808084e",	x"081307d1",	x"03726030",	
					x"07dd07b5",	x"07b607dc",	x"07d907ce",	x"07c707e4",	
					x"07d1082c",	x"07fa07ff",	x"080307f7",	x"07f207f2",	
					x"07f10821",	x"080b084d",	x"080f0815",	x"08090837",	
					x"0812082b",	x"084f083b",	x"080c0822",	x"07f70804",	
					x"07ea081f",	x"081b0826",	x"0808083a",	x"08430855",	
					x"082d0863",	x"084e086c",	x"083c085c",	x"08120847",	
					x"0807086b",	x"0854086b",	x"084a0881",	x"085d088b",	
					x"084608c0",	x"085c088b",	x"086b0891",	x"0867082f",	
					x"03727030",	x"081e07f4",	x"07de080d",	x"07c8080d",	
					x"07ed07ff",	x"082b0833",	x"0818088c",	x"087d0870",	
					x"08650842",	x"085408bf",	x"084b0886",	x"088d0885",	
					x"087508e5",	x"089c08bb",	x"089408ae",	x"08a30878",	
					x"089d086f",	x"087c08bf",	x"08b508ea",	x"08b208dd",	
					x"08b208f9",	x"08b608e3",	x"08c608c9",	x"089f08cd",	
					x"08a80894",	x"08b308fc",	x"08ff0909",	x"08f008e8",	
					x"090208fe",	x"08fc08fb",	x"08fc093c",	x"090b092c",	
					x"09010708",	x"000a0004",	x"9b18b16c",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"13730030",	x"071106b8",	x"06cc06f8",	
					x"06f606dd",	x"06e606fa",	x"06ff0713",	x"07070717",	
					x"0722071a",	x"072706e9",	x"06ec06ce",	x"070e0724",	
					x"07250718",	x"070d071c",	x"07470727",	x"07380734",	
					x"073c0720",	x"073b06d9",	x"06f506f0",	x"07180744",	
					x"07130721",	x"0738071f",	x"071a071e",	x"073a0726",	
					x"0713071e",	x"072d06bc",	x"06de0723",	x"07380738",	
					x"07300739",	x"070c071c",	x"07240735",	x"07130752",	
					x"07290710",	x"070506eb",	x"13731030",	x"06fa06b7",	
					x"06c306d2",	x"06d306c7",	x"06e906f7",	x"06ee0713",	
					x"070d0706",	x"071c0721",	x"07140716",	x"072c0723",	
					x"071e0712",	x"07300718",	x"07460715",	x"07360713",	
					x"0724071f",	x"071f071d",	x"072206b8",	x"06de06fc",	
					x"07130708",	x"071d071b",	x"07230721",	x"0717071b",	
					x"071806fd",	x"06ff06ff",	x"070006f8",	x"06d70706",	
					x"070d0721",	x"07230737",	x"07210714",	x"0735073d",	
					x"07370744",	x"0731074c",	x"073a06ca",	x"13732030",	
					x"06ca06dc",	x"06e706d6",	x"06dd06dc",	x"06d306cd",	
					x"06c806d4",	x"06f606f4",	x"071906de",	x"06ff06c3",	
					x"06ff06cc",	x"06f606d7",	x"07170712",	x"072906e3",	
					x"0705070c",	x"0708070f",	x"070d070c",	x"070606b8",	
					x"06cc06df",	x"06f206fb",	x"06f40714",	x"07310714",	
					x"0708070c",	x"06f90702",	x"07000715",	x"070206d4",	
					x"06d50704",	x"07110716",	x"0707071f",	x"0707071c",	
					x"07240722",	x"072f0722",	x"0722070d",	x"06fc06bf",	
					x"13733030",	x"06b306b1",	x"069306c7",	x"06e006ac",	
					x"06b106e1",	x"06e006e5",	x"06ea06f2",	x"06ec06ec",	
					x"06e806c2",	x"06e606ee",	x"06e306f5",	x"070506f9",	
					x"06ee06f0",	x"06e706ef",	x"06f706e5",	x"06f206dc",	
					x"06d806b3",	x"06b406eb",	x"06e106f9",	x"06f406fd",	
					x"07040712",	x"070c0724",	x"0721071b",	x"07160718",	
					x"071206e3",	x"06f30709",	x"07010720",	x"07090718",	
					x"07020728",	x"07090732",	x"071f0735",	x"070d0734",	
					x"06ff06a6",	x"000a0004",	x"54aa200f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"13744030",	x"06b506ae",	x"06b606db",	
					x"06bd06df",	x"06ea06ea",	x"06e906e3",	x"06df070b",	
					x"070b0714",	x"071306df",	x"06e10726",	x"07260727",	
					x"07360731",	x"072c072a",	x"0721072f",	x"073a0739",	
					x"0729072c",	x"07350704",	x"06ff0722",	x"072b0721",	
					x"07330744",	x"0764074b",	x"07460743",	x"0755074b",	
					x"074d072a",	x"072a0713",	x"0735074a",	x"07510759",	
					x"075f074f",	x"07580761",	x"07640760",	x"07630776",	
					x"075e0777",	x"0755071f",	x"13745030",	x"07260725",	
					x"071b0738",	x"07140703",	x"07260732",	x"07240737",	
					x"072c0750",	x"073d0764",	x"075c0715",	x"0732074e",	
					x"074a078d",	x"07660766",	x"075b075b",	x"07540756",	
					x"0750074d",	x"074c075e",	x"075a0727",	x"07080754",	
					x"07490767",	x"074b077d",	x"07750797",	x"076d0787",	
					x"076b0782",	x"075c077d",	x"07300761",	x"0758077e",	
					x"076d0792",	x"076d079c",	x"078b079b",	x"076a07aa",	
					x"079007a8",	x"078f07a0",	x"07760716",	x"13746030",	
					x"070d0739",	x"07180732",	x"07210713",	x"06fa0761",	
					x"071f075b",	x"0744075e",	x"0748074f",	x"0726076a",	
					x"07570769",	x"07820795",	x"07850784",	x"07950791",	
					x"07800796",	x"079307a8",	x"078007b0",	x"07870771",	
					x"075e07a1",	x"079e07aa",	x"079307b3",	x"07a507b4",	
					x"07a207d1",	x"079407bb",	x"079c07c6",	x"07c807a3",	
					x"07b707cd",	x"07c707d3",	x"07a707ed",	x"07c507fd",	
					x"07d007fe",	x"07c9080f",	x"07e307d4",	x"07ac0794",	
					x"13747030",	x"078a076e",	x"077207d2",	x"0762077f",	
					x"077007c0",	x"07a907de",	x"079707cf",	x"07c907df",	
					x"07df07cf",	x"07ba0812",	x"07d8080c",	x"07eb0809",	
					x"08150825",	x"0817081b",	x"0827082c",	x"081407f3",	
					x"07eb0804",	x"07df0814",	x"08230834",	x"081a084d",	
					x"083d0840",	x"082b0843",	x"08250846",	x"082c0838",	
					x"084e080f",	x"08310858",	x"08550854",	x"08500889",	
					x"085f0887",	x"08750884",	x"085e088e",	x"08670870",	
					x"08440776",	x"000a0004",	x"90d966ec",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"23750030",	x"079c0763",	x"076c0771",	
					x"076e0764",	x"07880795",	x"0798079e",	x"07b907d4",	
					x"07ca07ad",	x"07b6078e",	x"079e079e",	x"07c507c4",	
					x"07c107d2",	x"07d507c2",	x"07d80791",	x"0792079c",	
					x"079007ab",	x"0787074c",	x"07620793",	x"07af0785",	
					x"07830798",	x"07be07a9",	x"07a807ad",	x"079707b3",	
					x"07d007cf",	x"07ad0749",	x"077607a4",	x"07af07a1",	
					x"07aa07ad",	x"079907ab",	x"079907a6",	x"07b807c6",	
					x"07bd07d2",	x"07b90753",	x"23751030",	x"0781074a",	
					x"07530750",	x"076307a4",	x"07ac0775",	x"078e0786",	
					x"077e0778",	x"07a10781",	x"07810784",	x"079807b5",	
					x"07aa07c5",	x"07a007a7",	x"079d078d",	x"079c0775",	
					x"07900774",	x"0792074d",	x"07940750",	x"0775076a",	
					x"078707ab",	x"07a8078b",	x"07af0797",	x"079a078c",	
					x"079b0798",	x"07900787",	x"07b6075e",	x"0793078b",	
					x"079f07ae",	x"07ac07b9",	x"07a7077e",	x"07b607a5",	
					x"07b107bb",	x"07ba07b4",	x"07b10756",	x"23752030",	
					x"078a0727",	x"0715073d",	x"075e074f",	x"07890784",	
					x"07950767",	x"07800768",	x"07810768",	x"07830756",	
					x"07800768",	x"078f0780",	x"0791079f",	x"078e0786",	
					x"07920761",	x"07830797",	x"0796077e",	x"07630756",	
					x"073a075a",	x"07680771",	x"07800779",	x"07860758",	
					x"076f077f",	x"07800779",	x"0775077a",	x"075f0762",	
					x"0762076f",	x"076f076a",	x"0783078e",	x"078b0774",	
					x"07860792",	x"07880794",	x"07720786",	x"075c0700",	
					x"23753030",	x"073c071b",	x"070e072c",	x"07110724",	
					x"07270739",	x"0748072e",	x"074d0741",	x"07480743",	
					x"072f0734",	x"0761074b",	x"0753076c",	x"0778076f",	
					x"076a0771",	x"0753075f",	x"07560755",	x"076a075c",	
					x"07430713",	x"07590751",	x"07580765",	x"07530764",	
					x"07450761",	x"076e0765",	x"07760784",	x"07650780",	
					x"077a0738",	x"0730077d",	x"07580763",	x"07510782",	
					x"077c078a",	x"0772079e",	x"0777078d",	x"077a07a1",	
					x"0783073a",	x"000a0004",	x"d3125d19",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"23764030",	x"07510738",	x"073c0758",	
					x"07490729",	x"072c0742",	x"07650754",	x"0761075b",	
					x"07530767",	x"07690755",	x"07690784",	x"078e078d",	
					x"07800779",	x"0787077f",	x"0789077c",	x"079a078a",	
					x"07950773",	x"077f077d",	x"078c0783",	x"0795078f",	
					x"07a8078e",	x"07a1078e",	x"07aa078f",	x"07c207ab",	
					x"07bc07a8",	x"07b60781",	x"07a30784",	x"079607a1",	
					x"07ba07ab",	x"07c207ee",	x"07c407cd",	x"07c707be",	
					x"07c107b4",	x"07bd0753",	x"23765030",	x"07900767",	
					x"07600778",	x"07630785",	x"077907a7",	x"07a707b1",	
					x"07b507c1",	x"07c007a0",	x"07c107c1",	x"07b707ce",	
					x"07ab07e0",	x"07d407de",	x"07de07c0",	x"07bf07d3",	
					x"07e307c4",	x"07b607dd",	x"07a607b3",	x"079c07c3",	
					x"07d307ec",	x"07cf07ed",	x"07dc07f3",	x"07cb07f0",	
					x"07d007e4",	x"07ce07e1",	x"07b607c1",	x"07b107f2",	
					x"07d407fe",	x"07ec07fd",	x"07ea084c",	x"07db082d",	
					x"07fe0817",	x"07ed0803",	x"07de0796",	x"23766030",	
					x"0783079b",	x"078e07a8",	x"079d0797",	x"07ae07ed",	
					x"07af07b9",	x"07a707b5",	x"07a607a7",	x"07c707b8",	
					x"07e10804",	x"07ea080b",	x"07f10800",	x"080b0813",	
					x"07ce0810",	x"07ee080e",	x"07fd0810",	x"07fa0803",	
					x"07ef0801",	x"0804080d",	x"07f60818",	x"080e081d",	
					x"081c0847",	x"081d0815",	x"0800082b",	x"08090811",	
					x"080e083e",	x"0828082d",	x"08170846",	x"083a0864",	
					x"08270860",	x"08400862",	x"08180853",	x"081807ee",	
					x"23767030",	x"07d107bc",	x"07a107dc",	x"07d807dc",	
					x"07ef0848",	x"07ee080b",	x"08150846",	x"083b0844",	
					x"081e0844",	x"08370869",	x"0857086f",	x"086a085d",	
					x"085c0867",	x"085a0876",	x"08720888",	x"08810851",	
					x"0854086a",	x"08590882",	x"088008b1",	x"08900888",	
					x"088a08a0",	x"087e08a5",	x"08b708e4",	x"08a508a6",	
					x"08aa0885",	x"08a208c4",	x"08c008cf",	x"08b108cb",	
					x"08c508f3",	x"08ce08f3",	x"08e508f5",	x"08dd08d7",	
					x"08d706c7",	x"000a0004",	x"06aa98f8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"33770030",	x"071b06b0",	x"06b006be",	
					x"06bb06c8",	x"06d906c3",	x"070206d4",	x"07060710",	
					x"071e06e1",	x"070306dd",	x"06da06da",	x"07170741",	
					x"074d06e4",	x"070706e7",	x"06fc06f4",	x"072306ea",	
					x"06e706b7",	x"06c7069e",	x"06d806d8",	x"06db06da",	
					x"070406da",	x"070006fa",	x"070d0710",	x"07380704",	
					x"06f306e3",	x"070006e7",	x"06f6071f",	x"073306f4",	
					x"070406f3",	x"06fa06e3",	x"070a06ec",	x"070d0713",	
					x"07250729",	x"071a068c",	x"33771030",	x"06a30697",	
					x"069d06cc",	x"06d30692",	x"06ad06dc",	x"06d3070c",	
					x"06fa06db",	x"06ea06da",	x"06e206c5",	x"06e206f6",	
					x"06f4070e",	x"07290711",	x"0711070e",	x"070f06f1",	
					x"06e606f1",	x"06e606bb",	x"06d206cb",	x"06e506c8",	
					x"06ee06d0",	x"070306d6",	x"06f106f5",	x"071406e6",	
					x"072a06ff",	x"06fa06ff",	x"06ef06cc",	x"06ca06ec",	
					x"06f406e7",	x"06eb06ee",	x"06f70705",	x"070e0706",	
					x"07100717",	x"06ee0739",	x"0734068b",	x"33772030",	
					x"06bf0693",	x"069906a2",	x"06c806ad",	x"06b806ab",	
					x"06c706c7",	x"06d906bf",	x"06e606ac",	x"06fb06c3",	
					x"06e706d8",	x"06ef06c7",	x"06f706d6",	x"06f406e5",	
					x"06e406d5",	x"06ee06d4",	x"06e706d2",	x"06ef0693",	
					x"06c406ed",	x"06e306e1",	x"06e406e9",	x"06e706e4",	
					x"06d806d9",	x"06cc06f5",	x"06da06bb",	x"06b806ab",	
					x"06c206e7",	x"06d106f4",	x"06ee06de",	x"06e806e1",	
					x"06f806f9",	x"06f506fd",	x"06ec0703",	x"0701069a",	
					x"33773030",	x"06ae0682",	x"069f068b",	x"069606a0",	
					x"069806b9",	x"069a069a",	x"06bb06bf",	x"06c006ab",	
					x"06b806a9",	x"06b806cf",	x"06db06dd",	x"06c506fa",	
					x"06e706df",	x"06ca06ce",	x"06bc06c8",	x"06be06c7",	
					x"06da069e",	x"06a106cd",	x"06d006d5",	x"06cf06de",	
					x"06d906ee",	x"06d706f4",	x"06e806e4",	x"06d606f6",	
					x"06f406bb",	x"06ab06bc",	x"06c80711",	x"06d206f2",	
					x"06cb06f4",	x"06d10712",	x"06e60713",	x"06fd070e",	
					x"06df06c1",	x"000a0004",	x"c44c0d04",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"33784030",	x"06b606ad",	x"068206c3",	
					x"06ab06d1",	x"06cd06c4",	x"06aa06be",	x"06d606b2",	
					x"06b706c9",	x"06d406cb",	x"06ce06e9",	x"06f106f3",	
					x"070806ef",	x"070406d9",	x"06e206f8",	x"06fd06eb",	
					x"06ff06e9",	x"06f906c1",	x"06d906fa",	x"06e406f9",	
					x"070f0716",	x"07200714",	x"07160723",	x"071b0711",	
					x"0719070b",	x"06fe06fe",	x"06fd0708",	x"0705070c",	
					x"07190735",	x"072d072e",	x"07270759",	x"07470746",	
					x"0742074f",	x"073106f8",	x"33785030",	x"070106fa",	
					x"06da06ed",	x"06d006e5",	x"06e706fc",	x"06f606f5",	
					x"06e906f5",	x"0703073c",	x"070b0705",	x"0712071b",	
					x"071e0746",	x"07330747",	x"073d0731",	x"0722072c",	
					x"0727072c",	x"07250726",	x"071506d1",	x"07060727",	
					x"07300740",	x"072b073d",	x"073f074d",	x"0731074f",	
					x"07250758",	x"072d074f",	x"073b0753",	x"0729076a",	
					x"072f075f",	x"07300764",	x"07410775",	x"07410778",	
					x"074a076a",	x"0746077c",	x"07610732",	x"33786030",	
					x"07280716",	x"06f4070a",	x"06f90714",	x"070b074b",	
					x"072f0730",	x"070f0720",	x"07130723",	x"071f0723",	
					x"06ef075f",	x"07620777",	x"07570767",	x"074a076d",	
					x"07570762",	x"07610778",	x"075f0769",	x"0769073d",	
					x"072a076a",	x"075b076d",	x"07700793",	x"077a077f",	
					x"07740774",	x"0777079d",	x"07890796",	x"07730774",	
					x"07790797",	x"077e0796",	x"07640799",	x"077607a9",	
					x"078007ae",	x"078507d9",	x"078d07b1",	x"0771076f",	
					x"33787030",	x"074c0762",	x"07570744",	x"07550744",	
					x"072d076e",	x"073d074d",	x"075c078a",	x"078a079e",	
					x"078f07aa",	x"07a307c1",	x"07c307d2",	x"07cf07cf",	
					x"07c807e0",	x"07b907dd",	x"07e107d6",	x"07a207d2",	
					x"07d007c3",	x"07ac07c3",	x"07cd07e2",	x"07d407fe",	
					x"07f707e4",	x"07f607f3",	x"07f2080b",	x"07fd0811",	
					x"081307d8",	x"07d8080e",	x"08040828",	x"07fd0811",	
					x"07dd085d",	x"07f8084a",	x"083b0843",	x"08220834",	
					x"081507a1",	x"000a0004",	x"f6ed4ce2",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"03790031",	x"07920745",	x"0793078a",	
					x"0744074d",	x"0748074f",	x"074c074f",	x"07550760",	
					x"07470767",	x"07760730",	x"07870792",	x"078e0796",	
					x"079f07a4",	x"07a10796",	x"07bb0795",	x"07b207b5",	
					x"0791077b",	x"07b40761",	x"07760775",	x"07a00780",	
					x"07a60794",	x"079c079b",	x"0799078d",	x"07960789",	
					x"07a1078a",	x"07aa0765",	x"078007a1",	x"07be07a6",	
					x"079c07b3",	x"07bb0795",	x"078f07b8",	x"07a707a2",	
					x"077f07a6",	x"079a0769",	x"03791031",	x"07950765",	
					x"07530753",	x"07520745",	x"072b0702",	x"0718071e",	
					x"07290712",	x"07200755",	x"0756073d",	x"0762076b",	
					x"07770781",	x"07970771",	x"07920775",	x"078b0774",	
					x"0780078b",	x"0782077f",	x"077b0751",	x"07640775",	
					x"078a077c",	x"0781078c",	x"077a0789",	x"07980770",	
					x"07710797",	x"079d078b",	x"079f0753",	x"0756078b",	
					x"0799077b",	x"079707b6",	x"07c307a5",	x"07a407cd",	
					x"07af07a6",	x"07a807a4",	x"07710731",	x"03792031",	
					x"07340764",	x"0761075c",	x"0748071a",	x"074606ef",	
					x"071f0722",	x"0714073c",	x"0729074d",	x"0777073c",	
					x"075e0770",	x"0781077a",	x"076f0776",	x"0789073a",	
					x"07610767",	x"07850749",	x"074f0742",	x"07500724",	
					x"075f0793",	x"0783075e",	x"075f076d",	x"076e075e",	
					x"07490751",	x"0772077a",	x"075e07a0",	x"078c0767",	
					x"076c076d",	x"076d0779",	x"07890765",	x"07660790",	
					x"075a0799",	x"0784078a",	x"076c078b",	x"07840715",	
					x"03793031",	x"07140729",	x"0728073d",	x"0721072c",	
					x"07070738",	x"0725071f",	x"06f90723",	x"072c0761",	
					x"07680748",	x"073e074f",	x"075b0760",	x"0745076c",	
					x"07500760",	x"07540770",	x"07630750",	x"073a0779",	
					x"07370740",	x"074f0788",	x"0783078d",	x"07870789",	
					x"077c078a",	x"07780788",	x"0773078d",	x"07870798",	
					x"076d0780",	x"075b07a8",	x"076a0784",	x"07620792",	
					x"0786079c",	x"0786079b",	x"078307a1",	x"075007ae",	
					x"07720771",	x"000a0004",	x"497c572f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"037a4031",	x"074d075d",	x"07520774",	
					x"073c073a",	x"07220773",	x"072e0746",	x"07530757",	
					x"07540759",	x"074b0779",	x"073f0793",	x"076507a4",	
					x"078407ba",	x"079b0798",	x"078b07ac",	x"07a107b7",	
					x"07a607b9",	x"079c0795",	x"079e07c1",	x"079f07ce",	
					x"07aa07c7",	x"07b307d6",	x"07b807d6",	x"07b107cb",	
					x"07c407d9",	x"07aa07e2",	x"07b707e4",	x"07d10818",	
					x"07e007f9",	x"07eb07fa",	x"07d00815",	x"07e707fc",	
					x"07cd07f4",	x"07c2079b",	x"037a5031",	x"077d079d",	
					x"07a40787",	x"076a0783",	x"077907a8",	x"07670791",	
					x"078e07ae",	x"079e07b6",	x"07a807ac",	x"07c607f0",	
					x"07d507df",	x"07d507f2",	x"07df07e5",	x"07d407f3",	
					x"07d207f7",	x"07cb0806",	x"07c707c2",	x"07a607f3",	
					x"07e007f4",	x"07bb07f8",	x"07c207ff",	x"07d80836",	
					x"07e4083c",	x"07dd0821",	x"07d007f4",	x"07ee083d",	
					x"07f40826",	x"07f20835",	x"08070837",	x"07e1082e",	
					x"08010839",	x"07ef081b",	x"07e80796",	x"037a6031",	
					x"078407c0",	x"07b107fc",	x"07a307a9",	x"076e07c1",	
					x"078d07b5",	x"07ad07ed",	x"079707ea",	x"07e307ec",	
					x"07c5081e",	x"07e60826",	x"07fa0812",	x"07f4081b",	
					x"0803084b",	x"07f9082d",	x"08250844",	x"07f1080a",	
					x"07e50829",	x"08200815",	x"0807083c",	x"080d0871",	
					x"083d0880",	x"08320846",	x"08110877",	x"08190819",	
					x"08050881",	x"08340877",	x"0825087e",	x"08450877",	
					x"081e0882",	x"082d086d",	x"084c086d",	x"0849082d",	
					x"037a7031",	x"082a080a",	x"07db07ff",	x"07ad0815",	
					x"07d4080e",	x"07e00833",	x"07e3085e",	x"07f50851",	
					x"08200851",	x"082d0892",	x"0850088d",	x"08840894",	
					x"08930897",	x"087c08bf",	x"087a08c5",	x"086208a5",	
					x"08700878",	x"087b08b2",	x"088908be",	x"089b08c1",	
					x"088b08d3",	x"089508f4",	x"08af08f3",	x"08a008de",	
					x"08a308bd",	x"08a308f1",	x"08cb092e",	x"08f6091f",	
					x"08e908ff",	x"08d10900",	x"08f00915",	x"08be08fd",	
					x"08e906db",	x"000a0004",	x"89f0abf8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"137b0031",	x"07000717",	x"06f20715",	
					x"06f306ed",	x"06d706e6",	x"06dc06e8",	x"06e106db",	
					x"06de06c4",	x"06cd06d6",	x"06d506fa",	x"070e0706",	
					x"07110708",	x"070206f5",	x"0728070a",	x"072e0714",	
					x"07290709",	x"071806d0",	x"071f06e2",	x"070c072e",	
					x"07090713",	x"072c0717",	x"070d0726",	x"071b0716",	
					x"06ff0702",	x"073006df",	x"06d906ff",	x"0714072f",	
					x"070d0725",	x"0720071f",	x"06e10722",	x"07160731",	
					x"071d06f6",	x"07110709",	x"137b1031",	x"06fd06f8",	
					x"06fa06da",	x"06ee06c1",	x"06d206b4",	x"069706c0",	
					x"06c106e2",	x"06cb06d1",	x"06bc06b9",	x"06d00701",	
					x"06e70710",	x"06fd06f2",	x"070406ed",	x"070506ff",	
					x"071c071a",	x"070606ec",	x"070a06db",	x"06fc06e9",	
					x"06e00720",	x"07220703",	x"07090703",	x"071106ef",	
					x"070706f3",	x"06fd06f0",	x"070006fc",	x"06ea070e",	
					x"070f0715",	x"0709071c",	x"071f0711",	x"07200728",	
					x"0718072a",	x"0724073c",	x"072206bf",	x"137b2031",	
					x"06ed06d3",	x"06e106e6",	x"06c906c7",	x"06cf06be",	
					x"06cc06ad",	x"06a406b8",	x"06c606cc",	x"06ec06a5",	
					x"06e606b9",	x"070306f8",	x"07060713",	x"070f0706",	
					x"06f606f3",	x"070906f3",	x"070406f2",	x"06f906b5",	
					x"06d406ef",	x"06f906e9",	x"06fc06fb",	x"070506f8",	
					x"06e706fd",	x"06eb071a",	x"06f80702",	x"071306eb",	
					x"06d806f8",	x"0715071f",	x"07130711",	x"07060712",	
					x"070e071f",	x"072a0728",	x"07200723",	x"06e906cf",	
					x"137b3031",	x"06c506c4",	x"069406b8",	x"06a606ca",	
					x"06d206cd",	x"06af06a2",	x"06ac06ad",	x"06a70699",	
					x"069e0690",	x"069106da",	x"06d60702",	x"06d10712",	
					x"06f3070e",	x"06e606ec",	x"06d506fa",	x"06e806ec",	
					x"06df06e0",	x"06dc06fb",	x"070106ff",	x"0703070a",	
					x"06ff0716",	x"071b0712",	x"06f2070e",	x"070f070e",	
					x"070406f4",	x"06e40707",	x"06e80729",	x"07090731",	
					x"07010750",	x"07090734",	x"070b072b",	x"0703071b",	
					x"06e806e3",	x"000a0004",	x"4c221af8",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"137c4031",	x"06d606ec",	x"06df06fb",	
					x"06e206ff",	x"06ef06ce",	x"06c106e5",	x"06c606e4",	
					x"06d006f2",	x"06d006f3",	x"06ed0718",	x"070e0715",	
					x"0718073c",	x"0728071a",	x"0723072b",	x"07370740",	
					x"072a0734",	x"072d071e",	x"071f0729",	x"072f0752",	
					x"07400757",	x"074e0756",	x"073e073b",	x"073e076e",	
					x"0753074d",	x"0740072d",	x"072b0772",	x"07730781",	
					x"075e0783",	x"07700780",	x"07630791",	x"076507a0",	
					x"076d0779",	x"072a0718",	x"137c5031",	x"07060728",	
					x"0726074f",	x"071b074d",	x"07070742",	x"0722074c",	
					x"07130752",	x"07180745",	x"073b072b",	x"0721076f",	
					x"074a0789",	x"074e0780",	x"074e0775",	x"07700774",	
					x"075c077a",	x"075b0773",	x"07560768",	x"075b078c",	
					x"07740792",	x"0765077d",	x"076d07aa",	x"074707b0",	
					x"078907a4",	x"077207a2",	x"075a0784",	x"075807ac",	
					x"079807ba",	x"076407c8",	x"079207a9",	x"076907b7",	
					x"07a207a9",	x"077f079b",	x"076d0729",	x"137c6031",	
					x"0710074d",	x"073a075b",	x"0735074b",	x"07100751",	
					x"07330737",	x"07040749",	x"06ff0764",	x"07250742",	
					x"072e0795",	x"076b078d",	x"074a079a",	x"079107cb",	
					x"079207b6",	x"078e07b1",	x"077507ce",	x"077a0794",	
					x"078d07bb",	x"079b07c6",	x"079b07cd",	x"07bf07d3",	
					x"07ae07db",	x"07a607e2",	x"07a907b3",	x"079b07ac",	
					x"078807ee",	x"07c60803",	x"07ab07f5",	x"07b90808",	
					x"07c00801",	x"07d40800",	x"07b607e1",	x"07a0078b",	
					x"137c7031",	x"077b07ac",	x"078107c3",	x"079907a5",	
					x"079c07c0",	x"077407c5",	x"078707a7",	x"0768079e",	
					x"079907b0",	x"07a7080b",	x"07d60813",	x"07c80822",	
					x"0821081e",	x"08080829",	x"0820085b",	x"080f0810",	
					x"0806081b",	x"07e70845",	x"0816085f",	x"0816084e",	
					x"08220841",	x"0825084b",	x"082e086a",	x"0846084e",	
					x"0835081a",	x"08330869",	x"083508b0",	x"0843088c",	
					x"0850087e",	x"084f08a5",	x"087408a5",	x"08760882",	
					x"084f076f",	x"000a0004",	x"8f1c6f64",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"237d0031",	x"079d0787",	x"07810786",	
					x"0760071f",	x"07610760",	x"075f075e",	x"075d0785",	
					x"07840762",	x"0781078b",	x"0797078a",	x"078a0782",	
					x"0785079d",	x"078d0787",	x"07890799",	x"077b0798",	
					x"07bb07b3",	x"078c0745",	x"07800785",	x"07880785",	
					x"076d079b",	x"07880786",	x"07ac07a9",	x"07aa07aa",	
					x"07c107c9",	x"07c2079b",	x"077d07a7",	x"07a007a3",	
					x"07b607ba",	x"07b70797",	x"078a07a7",	x"079207b6",	
					x"078c07bf",	x"07a70773",	x"237d1031",	x"07780759",	
					x"074f073d",	x"074b075e",	x"074d071c",	x"07500754",	
					x"07390796",	x"077c076b",	x"077d075f",	x"076807af",	
					x"079f07a7",	x"078707a0",	x"07be0771",	x"0789077b",	
					x"07a10794",	x"07a10771",	x"078d0770",	x"0795077c",	
					x"0784077e",	x"07790771",	x"0793077a",	x"0788076c",	
					x"079207a2",	x"07920799",	x"07a30764",	x"078c077c",	
					x"07b707c1",	x"07d107a5",	x"079007ae",	x"07c007a9",	
					x"07b107b2",	x"079607ae",	x"079b0745",	x"237d2031",	
					x"07590759",	x"075e0728",	x"0738075e",	x"073e074c",	
					x"072b0749",	x"0747073c",	x"07620776",	x"077d0712",	
					x"07460779",	x"079a077c",	x"077c0769",	x"0763074e",	
					x"07690782",	x"078d0780",	x"0772077c",	x"0769074d",	
					x"075a0761",	x"075c0790",	x"0788077f",	x"07760762",	
					x"07660779",	x"07a50780",	x"077c0788",	x"076f077e",	
					x"076a07a5",	x"0770077d",	x"077a07a2",	x"0783077a",	
					x"0784078b",	x"07780790",	x"07880796",	x"076f071d",	
					x"237d3031",	x"072e0734",	x"0721074a",	x"07210724",	
					x"071e0724",	x"06fe071a",	x"07250741",	x"071e072f",	
					x"0720070f",	x"073b0777",	x"076d076e",	x"07640764",	
					x"07540766",	x"07430773",	x"074f0777",	x"0772077d",	
					x"076f073f",	x"07630766",	x"0784075a",	x"07560768",	
					x"0761078a",	x"07680794",	x"077f078f",	x"076c0793",	
					x"07770772",	x"074d07bd",	x"077f0799",	x"077e0797",	
					x"07710796",	x"077707a9",	x"077b0798",	x"078407aa",	
					x"0777073d",	x"000a0004",	x"cd435c0f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"237e4031",	x"07540763",	x"0714074f",	
					x"073b0753",	x"07540741",	x"073f075b",	x"076d076c",	
					x"07570764",	x"07570763",	x"076d079c",	x"077b078a",	
					x"077e078a",	x"077e0793",	x"07810792",	x"079807d0",	
					x"079807a3",	x"0787079e",	x"07ac07af",	x"07ae07a9",	
					x"07ca07d1",	x"07b007be",	x"07ba07c1",	x"07b007c8",	
					x"07c407e7",	x"07d707c0",	x"07c807eb",	x"07c507d5",	
					x"07cb07d8",	x"07df07c8",	x"07cc07eb",	x"07d007d3",	
					x"07c407db",	x"07df077c",	x"237e5031",	x"07780791",	
					x"07890798",	x"075d0797",	x"079007c6",	x"077b07b7",	
					x"077f07ba",	x"07a107ce",	x"079a07a1",	x"079107e5",	
					x"07cc07f3",	x"07cd07e4",	x"07d3080b",	x"07cf07ef",	
					x"07da080d",	x"07dc07f9",	x"07d207f5",	x"07a807ef",	
					x"07b1080e",	x"07b6080e",	x"07ef0822",	x"07e7081c",	
					x"07f30827",	x"07fe0827",	x"080907fd",	x"07e30839",	
					x"07da082f",	x"07e7082a",	x"07f10831",	x"07e5083f",	
					x"08130835",	x"080b0821",	x"07e40795",	x"237e6031",	
					x"078307a3",	x"0788079f",	x"077607bb",	x"077d07e3",	
					x"079307b1",	x"077f07d5",	x"07ba07d6",	x"07b507cd",	
					x"07c707fc",	x"07f40818",	x"07d70825",	x"07e8084e",	
					x"07e6083d",	x"07ea0822",	x"07f9083d",	x"07e70837",	
					x"07f90820",	x"08100841",	x"0811084f",	x"081d0853",	
					x"08210897",	x"0829088e",	x"08370851",	x"082a0861",	
					x"0832085d",	x"08380842",	x"082f085f",	x"0823086a",	
					x"080c0868",	x"0834086f",	x"082d0857",	x"083807fc",	
					x"237e7031",	x"07d90819",	x"08090825",	x"07cb0842",	
					x"07d10840",	x"07f7082c",	x"08120862",	x"081c0883",	
					x"082f0841",	x"083c0882",	x"086f089b",	x"088e0898",	
					x"086a08a4",	x"0868089f",	x"088008b1",	x"089408ad",	
					x"08770888",	x"086a08ba",	x"089e08ce",	x"089208c0",	
					x"089308d1",	x"089508d2",	x"08c708d6",	x"08cc08ce",	
					x"08d308c8",	x"08c408e4",	x"08ca08d6",	x"08bc08ea",	
					x"08cf08fb",	x"08a60906",	x"08db0910",	x"08df08f3",	
					x"08e50702",	x"000a0004",	x"0a50aa3e",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"337f0031",	x"071306b0",	x"06a006cd",	
					x"06b706a3",	x"068a06b6",	x"06be06ac",	x"06c506c8",	
					x"06c306ac",	x"06b806a8",	x"06b406f3",	x"070106e7",	
					x"071a06e3",	x"071a0700",	x"06f706ea",	x"07200701",	
					x"071506ef",	x"06ea06bf",	x"06fb06ec",	x"06f2070a",	
					x"07160703",	x"070506e9",	x"070006f5",	x"06fb0700",	
					x"071206f1",	x"073406dc",	x"070206eb",	x"0705070b",	
					x"0710070e",	x"070806e4",	x"070f06e6",	x"06f2072a",	
					x"0710070d",	x"070406b9",	x"337f1031",	x"06a506ce",	
					x"06bf06b1",	x"06a7069f",	x"06a006a6",	x"06a106a2",	
					x"06af0699",	x"06c806eb",	x"06e4069c",	x"06b906cb",	
					x"06e506f0",	x"06e006e9",	x"06dc06dc",	x"06d206db",	
					x"06f006f0",	x"06df06c3",	x"06be06c0",	x"06db06f0",	
					x"070a06d7",	x"06f406d9",	x"06fd06e5",	x"06fd06da",	
					x"06fc071b",	x"07040717",	x"070b06ca",	x"06d806fd",	
					x"07080704",	x"06fa06ef",	x"070d0710",	x"070806fb",	
					x"06f7072c",	x"070d0719",	x"070906bd",	x"337f2031",	
					x"06bc06c5",	x"06cf06aa",	x"06a506c7",	x"06ae0690",	
					x"0694069c",	x"06a306af",	x"06c706b5",	x"06dd06ad",	
					x"06c306db",	x"06e606db",	x"06ec06dd",	x"06fa06c8",	
					x"06de06dd",	x"06ef06e8",	x"06e606f0",	x"06e306b5",	
					x"06c306ea",	x"06e10703",	x"06e806e0",	x"06d806da",	
					x"06d506d2",	x"06d006e9",	x"06f006d8",	x"06c706d0",	
					x"06e5070c",	x"070006f0",	x"06e706f0",	x"06be06f2",	
					x"06d506ef",	x"06e706fb",	x"06db06fa",	x"06e306bb",	
					x"337f3031",	x"06b2068f",	x"0693068c",	x"066b06a8",	
					x"067f06bf",	x"066f0676",	x"068006c0",	x"06b0069d",	
					x"068c06a2",	x"06ae06ba",	x"06b506d7",	x"06a806e0",	
					x"06d006e0",	x"06d106dc",	x"06c306d5",	x"06c706dc",	
					x"06d506cc",	x"06ac06db",	x"06d006e7",	x"06dd06f8",	
					x"06eb06fd",	x"06e306e6",	x"06f50714",	x"06ef0709",	
					x"06d106f5",	x"06d80701",	x"06e706fc",	x"06dd06ff",	
					x"06ee070d",	x"06eb071c",	x"06cb0709",	x"06ee070c",	
					x"06e506b4",	x"000a0004",	x"bf890d9f",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"00c0ffee",	
					x"0000d125",	x"33804031",	x"06a006b9",	x"067a06cd",	
					x"068106d5",	x"069e06db",	x"069906cd",	x"06a806f4",	
					x"06ba06c3",	x"06a706cf",	x"06cf0704",	x"06e80712",	
					x"070206ff",	x"06fb06f7",	x"06e6071c",	x"0703070f",	
					x"070a0710",	x"071506f5",	x"06f80732",	x"071b0709",	
					x"07080725",	x"07320726",	x"07280735",	x"071b073c",	
					x"0710074c",	x"07280735",	x"071c0732",	x"07140731",	
					x"071b073e",	x"071d073e",	x"072c075b",	x"0745077a",	
					x"0740074a",	x"071d06e8",	x"33805031",	x"06f6072e",	
					x"06dd06fc",	x"06b306fc",	x"06c906f9",	x"06d806f5",	
					x"06d20722",	x"07100712",	x"06ee0709",	x"07010739",	
					x"0720073d",	x"07360744",	x"0739073b",	x"0730075d",	
					x"07450742",	x"07280742",	x"07400727",	x"0720074a",	
					x"07390756",	x"073a075d",	x"07580774",	x"0750079b",	
					x"07400784",	x"07430779",	x"07400762",	x"07430799",	
					x"07500784",	x"074d077d",	x"074b076e",	x"07410782",	
					x"075607c5",	x"074e0777",	x"07620709",	x"33806031",	
					x"06fd071d",	x"06f40717",	x"06e3070a",	x"06de0719",	
					x"06f40711",	x"070d073d",	x"0712073c",	x"0741073f",	
					x"072c075f",	x"073f0790",	x"075b0777",	x"0754077b",	
					x"0769076e",	x"0772079c",	x"07700798",	x"075f0779",	
					x"07570779",	x"0783078b",	x"077b0794",	x"078f07b4",	
					x"076a0789",	x"077e07a2",	x"078007c8",	x"079007a2",	
					x"076e07d4",	x"079a07c8",	x"078a07d0",	x"079707d7",	
					x"078f07dc",	x"07ac07d8",	x"07a407b3",	x"077f074c",	
					x"33807031",	x"07540773",	x"075b079a",	x"07340767",	
					x"071e07bf",	x"0724079f",	x"076107a4",	x"07630791",	
					x"0768078c",	x"076d07ee",	x"07af07f6",	x"07c207e2",	
					x"07ba07fa",	x"07a707ec",	x"07d407f3",	x"07b107f2",	
					x"07cc07f2",	x"07cb080f",	x"07f8081f",	x"07cf07fd",	
					x"07f70808",	x"08000811",	x"07fd0823",	x"07fc081a",	
					x"07f60808",	x"0802083e",	x"081a0816",	x"07f30865",	
					x"08180856",	x"0806085e",	x"0820085e",	x"082e084c",	
					x"08140742",	x"000a0004",	x"f86e5936",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"ce11b10c",	
					x"0000d125",	x"00810000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"99999999",	x"99999999",	
					x"99999999",	x"000a0004",	x"1e89bcc5",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"000ab0de",	
					x"0000d125",	x"00820000",	x"03e803e8",	x"03e803e8",	
					x"03e803e8",	x"03e803e8",	x"03e803e8",	x"03e803e8",	
					x"03e803e8",	x"03e803e8",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"079e079e",	x"079e079e",	
					x"079e079e",	x"079e079e",	x"051e051e",	x"051e051e",	
					x"051e051e",	x"051e051e",	x"051e051e",	x"051e051e",	
					x"051e051e",	x"051e051e",	x"0c9e0c9e",	x"0c9e0c9e",	
					x"0c9e0c9e",	x"0c9e0c9e",	x"0c9e0c9e",	x"0c9e0c9e",	
					x"0c9e0c9e",	x"0c9e0c9e",	x"042e042e",	x"042e042e",	
					x"042e042e",	x"042e042e",	x"042e042e",	x"042e042e",	
					x"042e042e",	x"042e042e",	x"044c044c",	x"044c044c",	
					x"044c044c",	x"044c044c",	x"044c044c",	x"044c044c",	
					x"044c044c",	x"044c044c",	x"06400640",	x"06400640",	
					x"06400640",	x"06400640",	x"06400640",	x"06400640",	
					x"06400640",	x"06400640",	x"044c044c",	x"044c044c",	
					x"044c044c",	x"044c044c",	x"044c044c",	x"044c044c",	
					x"044c044c",	x"044c044c",	x"09130883",	x"09a909c8",	
					x"09ea085a",	x"08de099d",	x"0a2f0e7a",	x"0c450c8b",	
					x"0c7c0afd",	x"09820e24",	x"03840384",	x"03840384",	
					x"03840384",	x"03840384",	x"03840384",	x"03840384",	
					x"03840384",	x"03840384",	x"0ce40ce4",	x"0ce40ce4",	
					x"0ce40ce4",	x"0ce40ce4",	x"0ce40ce4",	x"0ce40ce4",	
					x"0ce40ce4",	x"0ce40ce4",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"0000050f",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"000a0004",	x"9200098d",	x"62504944",	
					x"00be11e2",	x"0000008c",	x"20111213",	x"000f00da",	
					x"0000d125",	x"00830000",	x"0000ffff",	x"0000079d",	
					x"0000079c",	x"0000079e",	x"0000079d",	x"000007a8",	
					x"0000079c",	x"0000079e",	x"000007a1",	x"0000079d",	
					x"0000079c",	x"0000079c",	x"0000079c",	x"0000079d",	
					x"0000079d",	x"0000079d",	x"00000799",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"00000000",	x"00000000",	x"00000000",	x"00000000",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"99999999",	x"99999999",	x"99999999",	
					x"99999999",	x"000a0004",	x"b6f0ec98",	x"62504944"	
				);
end data32_pkg;