x"00be11e2",	x"0000008c",	x"20111213",	x"0000eada",	
x"0000d125",	x"00000000",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"99999999",	x"99999999",	x"99999999",	
x"99999999",	x"000a0004",	x"1cc4c313",	x"62504944"
