library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package data16_pkg is

	type ram_type is array (0 to 132*(2*140)-1) of std_logic_vector(15 downto 0);
	constant data16 : ram_type :=(
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"eada",	x"0000",	
												x"d125",	x"0000",	x"0000",	x"0000",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"0004",	x"000a",	
												x"c313",	x"1cc4",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"0001",	
												x"06a5",	x"06d0",	x"06a5",	x"069f",	
												x"06a4",	x"068c",	x"069e",	x"06a4",	
												x"06ae",	x"0694",	x"06af",	x"068b",	
												x"0705",	x"06d4",	x"06ad",	x"06cf",	
												x"06d1",	x"06d3",	x"06d9",	x"06f2",	
												x"06f8",	x"06e6",	x"06b4",	x"06eb",	
												x"06e6",	x"06c8",	x"0703",	x"070c",	
												x"06f2",	x"0708",	x"06b3",	x"06f6",	
												x"06c3",	x"06c2",	x"06ee",	x"06e2",	
												x"06d9",	x"0702",	x"06e5",	x"06d9",	
												x"06c2",	x"06d4",	x"06f8",	x"06de",	
												x"06e1",	x"06fc",	x"06a2",	x"06e5",	
												x"06e1",	x"06c7",	x"06de",	x"06d8",	
												x"06f1",	x"06d3",	x"071f",	x"06f6",	
												x"06bc",	x"06c9",	x"06f3",	x"06e1",	
												x"0706",	x"06cd",	x"067b",	x"06e4",	
												x"102e",	x"0001",	x"0685",	x"069e",	
												x"06b1",	x"069f",	x"0667",	x"06a2",	
												x"067a",	x"068d",	x"06b3",	x"068b",	
												x"06b0",	x"06b2",	x"0696",	x"06b0",	
												x"069c",	x"06b6",	x"06dd",	x"068d",	
												x"06d7",	x"06e8",	x"06be",	x"06ce",	
												x"06c5",	x"06dd",	x"06ae",	x"06cd",	
												x"06cb",	x"06bd",	x"06c9",	x"06be",	
												x"0678",	x"06d7",	x"06d7",	x"06c6",	
												x"06d7",	x"06df",	x"06ce",	x"06d6",	
												x"06ac",	x"06f4",	x"06ba",	x"06d2",	
												x"06dc",	x"06db",	x"06bf",	x"06d2",	
												x"06b4",	x"06c7",	x"06fb",	x"06d9",	
												x"06f8",	x"06e5",	x"06fe",	x"06eb",	
												x"06e9",	x"0706",	x"0701",	x"06f7",	
												x"0701",	x"0711",	x"06ec",	x"0706",	
												x"06aa",	x"06eb",	x"202e",	x"0001",	
												x"0695",	x"067e",	x"0692",	x"068c",	
												x"0676",	x"069c",	x"0691",	x"0680",	
												x"06a7",	x"0696",	x"06a3",	x"06c1",	
												x"06b2",	x"06a3",	x"069a",	x"06af",	
												x"06c5",	x"06c1",	x"06b6",	x"06d5",	
												x"06bf",	x"06d2",	x"06c0",	x"06d5",	
												x"06e7",	x"06c3",	x"06bc",	x"06ef",	
												x"06ac",	x"06b1",	x"068e",	x"06ac",	
												x"06aa",	x"068d",	x"06c6",	x"06a1",	
												x"06bd",	x"06be",	x"06c5",	x"06c3",	
												x"06d1",	x"06cd",	x"06cb",	x"06d8",	
												x"06c7",	x"06c8",	x"06ae",	x"06bc",	
												x"06d1",	x"06cd",	x"06d4",	x"06cc",	
												x"06e9",	x"06d3",	x"06ea",	x"06eb",	
												x"06ce",	x"06f1",	x"06c5",	x"06d4",	
												x"06dc",	x"069d",	x"065c",	x"06d2",	
												x"302e",	x"0001",	x"0668",	x"0651",	
												x"068a",	x"0672",	x"0694",	x"0688",	
												x"0674",	x"066f",	x"068c",	x"065d",	
												x"06b0",	x"069b",	x"06a0",	x"06a3",	
												x"067f",	x"0699",	x"06c7",	x"067d",	
												x"06c4",	x"06be",	x"06ca",	x"06be",	
												x"06dc",	x"06c3",	x"06db",	x"06b1",	
												x"06c5",	x"06ad",	x"06bf",	x"06c4",	
												x"0685",	x"06b7",	x"06be",	x"069c",	
												x"06c3",	x"06c0",	x"06c1",	x"06c3",	
												x"06cb",	x"06c6",	x"06c7",	x"06b5",	
												x"06cf",	x"06bb",	x"06d5",	x"06bd",	
												x"06bc",	x"06bc",	x"06ef",	x"06b5",	
												x"06da",	x"06bc",	x"06f4",	x"06c3",	
												x"06ec",	x"06db",	x"0705",	x"06cd",	
												x"06f6",	x"06cf",	x"06f2",	x"06c4",	
												x"069d",	x"06cf",	x"0004",	x"000a",	
												x"00b0",	x"e549",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"0002",	
												x"06b0",	x"067f",	x"0693",	x"0699",	
												x"06a9",	x"0689",	x"06d9",	x"0697",	
												x"06c5",	x"06a6",	x"06ee",	x"06ad",	
												x"06eb",	x"06d5",	x"06ae",	x"06cc",	
												x"06eb",	x"06c9",	x"06e4",	x"06ed",	
												x"06e2",	x"06ca",	x"06fb",	x"06e5",	
												x"06e4",	x"06d6",	x"06e8",	x"06ee",	
												x"06f3",	x"0704",	x"06ce",	x"06de",	
												x"070f",	x"06e0",	x"06fc",	x"0717",	
												x"0702",	x"06ed",	x"0710",	x"0700",	
												x"071b",	x"06f8",	x"06fe",	x"070a",	
												x"06f9",	x"06f9",	x"06fa",	x"06e8",	
												x"0713",	x"0705",	x"071f",	x"0706",	
												x"0721",	x"0712",	x"072d",	x"072a",	
												x"073f",	x"06ff",	x"0733",	x"071e",	
												x"072f",	x"06f6",	x"06e3",	x"070f",	
												x"502e",	x"0002",	x"06d1",	x"06ae",	
												x"06d9",	x"06a2",	x"06db",	x"06ad",	
												x"06ec",	x"06c6",	x"070d",	x"06e8",	
												x"070e",	x"06f5",	x"0710",	x"06f8",	
												x"0723",	x"06f7",	x"072c",	x"0704",	
												x"073c",	x"0720",	x"072a",	x"0730",	
												x"0733",	x"071b",	x"0724",	x"06ea",	
												x"073f",	x"072a",	x"0731",	x"06ee",	
												x"070b",	x"0702",	x"072d",	x"0712",	
												x"0749",	x"0713",	x"073d",	x"0717",	
												x"0739",	x"0723",	x"0740",	x"071f",	
												x"0745",	x"0718",	x"0755",	x"071d",	
												x"073d",	x"0716",	x"074a",	x"0709",	
												x"0770",	x"0735",	x"075d",	x"0739",	
												x"0774",	x"0721",	x"0763",	x"072d",	
												x"076f",	x"0731",	x"0752",	x"0726",	
												x"0700",	x"070b",	x"602e",	x"0002",	
												x"0715",	x"06c4",	x"0713",	x"06dd",	
												x"070a",	x"06d5",	x"072d",	x"06fa",	
												x"0724",	x"06ea",	x"0715",	x"06f6",	
												x"072c",	x"06f0",	x"072c",	x"06fd",	
												x"0743",	x"0708",	x"0741",	x"0734",	
												x"073a",	x"072e",	x"0768",	x"073c",	
												x"0757",	x"0736",	x"076b",	x"075f",	
												x"076d",	x"074f",	x"0743",	x"073d",	
												x"0774",	x"0729",	x"0763",	x"075b",	
												x"0773",	x"0758",	x"0770",	x"075a",	
												x"075d",	x"0753",	x"0776",	x"0753",	
												x"077f",	x"0752",	x"0756",	x"076f",	
												x"0782",	x"0751",	x"0781",	x"0761",	
												x"0787",	x"0742",	x"079a",	x"0760",	
												x"07a6",	x"074f",	x"0782",	x"0751",	
												x"078f",	x"075a",	x"0754",	x"075d",	
												x"702e",	x"0002",	x"075b",	x"071f",	
												x"0731",	x"071a",	x"072d",	x"06e2",	
												x"077a",	x"0718",	x"0765",	x"0729",	
												x"078b",	x"0734",	x"076d",	x"075e",	
												x"0752",	x"0753",	x"077f",	x"073b",	
												x"07ae",	x"0793",	x"07a6",	x"0788",	
												x"07b7",	x"0779",	x"07a9",	x"075b",	
												x"07c7",	x"07a2",	x"07b3",	x"0779",	
												x"07ae",	x"0781",	x"07be",	x"0782",	
												x"07c5",	x"078a",	x"07cf",	x"07a3",	
												x"07ea",	x"078a",	x"07d3",	x"07a0",	
												x"07c9",	x"07b2",	x"07be",	x"0799",	
												x"07bb",	x"07c0",	x"07ef",	x"07af",	
												x"0811",	x"07dd",	x"07fd",	x"07d6",	
												x"0800",	x"07e5",	x"0819",	x"07c1",	
												x"0821",	x"07e3",	x"0810",	x"0802",	
												x"0630",	x"07ea",	x"0004",	x"000a",	
												x"43fe",	x"185f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"1003",	
												x"0644",	x"0633",	x"064a",	x"0661",	
												x"063b",	x"0665",	x"064f",	x"0651",	
												x"0693",	x"0651",	x"0686",	x"069a",	
												x"068e",	x"066f",	x"0676",	x"068e",	
												x"066b",	x"0674",	x"0689",	x"0687",	
												x"067c",	x"0690",	x"06b2",	x"06a6",	
												x"06b1",	x"068e",	x"0692",	x"06cd",	
												x"068f",	x"06a3",	x"0660",	x"068c",	
												x"069d",	x"0669",	x"069b",	x"06a3",	
												x"0681",	x"0677",	x"0690",	x"0692",	
												x"06a9",	x"0692",	x"06bc",	x"06a6",	
												x"0689",	x"06b5",	x"066c",	x"06af",	
												x"06a6",	x"06a0",	x"06b8",	x"06a3",	
												x"06ba",	x"06b5",	x"06ad",	x"06aa",	
												x"06a2",	x"0696",	x"06a9",	x"068b",	
												x"06c7",	x"068b",	x"0603",	x"068c",	
												x"102e",	x"1003",	x"0624",	x"060c",	
												x"066c",	x"062a",	x"0645",	x"065a",	
												x"066f",	x"065f",	x"065b",	x"0662",	
												x"0663",	x"0668",	x"066a",	x"0666",	
												x"0652",	x"066b",	x"0684",	x"066a",	
												x"0690",	x"06a2",	x"068e",	x"0692",	
												x"068f",	x"0698",	x"067d",	x"0694",	
												x"068b",	x"0694",	x"0696",	x"0688",	
												x"0662",	x"06aa",	x"0661",	x"067b",	
												x"0683",	x"068b",	x"06ad",	x"067f",	
												x"065f",	x"06b0",	x"0676",	x"0656",	
												x"0693",	x"067b",	x"0675",	x"0695",	
												x"065a",	x"0685",	x"068f",	x"067c",	
												x"06a4",	x"0691",	x"06b7",	x"06a1",	
												x"06a3",	x"0699",	x"06a2",	x"069d",	
												x"06a5",	x"069a",	x"069b",	x"068f",	
												x"0631",	x"0685",	x"202e",	x"1003",	
												x"0626",	x"063e",	x"066c",	x"0631",	
												x"064b",	x"062a",	x"064a",	x"0652",	
												x"0656",	x"0664",	x"0651",	x"0671",	
												x"0655",	x"064f",	x"063c",	x"0670",	
												x"0660",	x"066f",	x"0645",	x"0678",	
												x"0666",	x"065c",	x"0673",	x"0670",	
												x"0680",	x"0678",	x"066b",	x"068e",	
												x"067b",	x"0691",	x"0628",	x"0668",	
												x"0661",	x"0653",	x"066d",	x"065a",	
												x"0673",	x"065c",	x"067e",	x"0682",	
												x"0698",	x"068d",	x"0699",	x"0684",	
												x"0691",	x"0680",	x"0662",	x"067e",	
												x"066d",	x"0685",	x"0672",	x"0684",	
												x"0684",	x"0678",	x"069b",	x"067a",	
												x"067d",	x"0684",	x"0688",	x"0682",	
												x"068a",	x"0677",	x"0635",	x"0667",	
												x"302e",	x"1003",	x"0644",	x"05ff",	
												x"0637",	x"062f",	x"0645",	x"0611",	
												x"064e",	x"0621",	x"0668",	x"064b",	
												x"0653",	x"0650",	x"0680",	x"0634",	
												x"0653",	x"0664",	x"0650",	x"063b",	
												x"0670",	x"066a",	x"0664",	x"065f",	
												x"0679",	x"065c",	x"0683",	x"066d",	
												x"066d",	x"0679",	x"0669",	x"0669",	
												x"0641",	x"064a",	x"0668",	x"0648",	
												x"067b",	x"066d",	x"0677",	x"0673",	
												x"067d",	x"067f",	x"0683",	x"067a",	
												x"067e",	x"0668",	x"067b",	x"0687",	
												x"066b",	x"066a",	x"0686",	x"0665",	
												x"0688",	x"0663",	x"06a3",	x"066e",	
												x"06a8",	x"0693",	x"06a8",	x"068c",	
												x"069a",	x"0694",	x"0693",	x"066b",	
												x"0626",	x"0673",	x"0004",	x"000a",	
												x"dae6",	x"feb5",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"1004",	
												x"064a",	x"060c",	x"0661",	x"0624",	
												x"065f",	x"0647",	x"067e",	x"064f",	
												x"0681",	x"0667",	x"067e",	x"0680",	
												x"0688",	x"0686",	x"067d",	x"067c",	
												x"0696",	x"066d",	x"068c",	x"067e",	
												x"0696",	x"0677",	x"0689",	x"0698",	
												x"06a8",	x"0690",	x"06a7",	x"06aa",	
												x"069a",	x"06a7",	x"0668",	x"06a3",	
												x"06aa",	x"0673",	x"06a5",	x"06ad",	
												x"06b3",	x"0694",	x"06cd",	x"06cb",	
												x"069c",	x"06ca",	x"06cd",	x"06a3",	
												x"06c6",	x"06b3",	x"069f",	x"06b0",	
												x"06c0",	x"06a7",	x"06e8",	x"06c3",	
												x"06d2",	x"06d9",	x"06dd",	x"06d2",	
												x"06ce",	x"06bd",	x"06d5",	x"06d0",	
												x"06cb",	x"06b6",	x"0697",	x"06bb",	
												x"502e",	x"1004",	x"067f",	x"0661",	
												x"0699",	x"0673",	x"0696",	x"0665",	
												x"06b6",	x"0699",	x"06bc",	x"067f",	
												x"06d7",	x"069c",	x"06bd",	x"06ba",	
												x"06c0",	x"06b6",	x"06dc",	x"069c",	
												x"06d8",	x"06d1",	x"06c2",	x"06bd",	
												x"06d3",	x"06cf",	x"06d9",	x"06b8",	
												x"06c7",	x"06d0",	x"06c3",	x"06b6",	
												x"0697",	x"06ae",	x"06d5",	x"068b",	
												x"06e1",	x"06b2",	x"06dd",	x"06d8",	
												x"06e7",	x"06ca",	x"06eb",	x"06ca",	
												x"06ed",	x"06cf",	x"06fd",	x"06df",	
												x"06c9",	x"06cd",	x"06df",	x"06ca",	
												x"070f",	x"06b7",	x"06ff",	x"06d9",	
												x"0700",	x"06e6",	x"06fe",	x"06d6",	
												x"0703",	x"06e1",	x"06f7",	x"06df",	
												x"0688",	x"06ec",	x"602e",	x"1004",	
												x"069d",	x"0654",	x"06ae",	x"0683",	
												x"06b7",	x"069b",	x"06c9",	x"0688",	
												x"06d5",	x"06b0",	x"06ce",	x"069f",	
												x"06c9",	x"06a2",	x"06b9",	x"06b1",	
												x"06d5",	x"069b",	x"06f6",	x"06c3",	
												x"0715",	x"06c7",	x"0712",	x"06fc",	
												x"070f",	x"06ea",	x"0701",	x"06db",	
												x"0710",	x"06c5",	x"06de",	x"06ef",	
												x"070f",	x"06ee",	x"0701",	x"070b",	
												x"0710",	x"06d8",	x"0714",	x"06e8",	
												x"0722",	x"06e9",	x"0710",	x"0724",	
												x"0714",	x"06ec",	x"0713",	x"0701",	
												x"0728",	x"06f5",	x"072b",	x"0704",	
												x"0731",	x"0703",	x"0730",	x"0705",	
												x"0747",	x"06e7",	x"073e",	x"0729",	
												x"071e",	x"0708",	x"06ba",	x"06fa",	
												x"702e",	x"1004",	x"06d5",	x"069e",	
												x"0702",	x"069d",	x"06e6",	x"06c4",	
												x"071e",	x"06c4",	x"06ee",	x"06db",	
												x"06e1",	x"06d9",	x"073a",	x"06de",	
												x"070d",	x"06d6",	x"0741",	x"070e",	
												x"0743",	x"071c",	x"0747",	x"071b",	
												x"077e",	x"0731",	x"074c",	x"0737",	
												x"074e",	x"074c",	x"0739",	x"0738",	
												x"073f",	x"0741",	x"0729",	x"071c",	
												x"0767",	x"074d",	x"076c",	x"0731",	
												x"0780",	x"0744",	x"0799",	x"0760",	
												x"0776",	x"0761",	x"0791",	x"0757",	
												x"0748",	x"076b",	x"0767",	x"072d",	
												x"077a",	x"0767",	x"07aa",	x"0785",	
												x"07c7",	x"077c",	x"079a",	x"0782",	
												x"07a4",	x"0786",	x"0782",	x"077f",	
												x"0712",	x"0776",	x"0004",	x"000a",	
												x"1739",	x"2e43",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"2005",	
												x"071e",	x"070c",	x"0712",	x"071b",	
												x"06ee",	x"06f7",	x"0740",	x"0710",	
												x"0754",	x"0734",	x"0745",	x"073d",	
												x"0729",	x"074d",	x"0719",	x"072d",	
												x"071d",	x"0747",	x"0751",	x"0738",	
												x"0764",	x"0750",	x"0797",	x"0795",	
												x"075f",	x"0787",	x"0787",	x"0765",	
												x"0745",	x"0790",	x"072b",	x"0757",	
												x"073c",	x"073f",	x"0750",	x"075c",	
												x"0746",	x"074c",	x"0784",	x"0767",	
												x"0742",	x"0765",	x"0765",	x"0762",	
												x"0769",	x"0778",	x"0738",	x"0772",	
												x"0759",	x"0752",	x"0761",	x"0746",	
												x"0763",	x"076d",	x"076f",	x"0780",	
												x"074d",	x"0762",	x"0765",	x"074c",	
												x"076a",	x"0756",	x"06e4",	x"0736",	
												x"102e",	x"2005",	x"06e5",	x"06e4",	
												x"06ff",	x"06cd",	x"072c",	x"06f7",	
												x"072f",	x"072d",	x"0701",	x"0755",	
												x"074c",	x"072c",	x"072c",	x"0738",	
												x"071e",	x"0743",	x"0751",	x"0744",	
												x"0741",	x"0741",	x"0759",	x"0759",	
												x"0795",	x"076d",	x"0740",	x"0772",	
												x"074e",	x"075d",	x"074f",	x"0754",	
												x"070e",	x"0742",	x"0739",	x"074b",	
												x"074c",	x"0747",	x"0737",	x"074b",	
												x"073c",	x"0739",	x"074b",	x"0727",	
												x"0795",	x"0772",	x"0763",	x"0772",	
												x"0730",	x"0768",	x"0753",	x"075a",	
												x"0743",	x"0756",	x"076f",	x"074f",	
												x"076d",	x"0768",	x"0762",	x"0765",	
												x"076a",	x"0762",	x"0755",	x"076d",	
												x"06f6",	x"0764",	x"202e",	x"2005",	
												x"06ed",	x"0703",	x"06d4",	x"06ed",	
												x"06d6",	x"06ea",	x"06f3",	x"06f8",	
												x"072e",	x"0709",	x"0721",	x"074d",	
												x"0726",	x"0726",	x"071b",	x"0750",	
												x"0711",	x"073d",	x"0721",	x"073f",	
												x"074d",	x"074f",	x"0757",	x"0752",	
												x"0762",	x"075e",	x"0749",	x"0769",	
												x"075b",	x"0747",	x"06d8",	x"074e",	
												x"0741",	x"0724",	x"074a",	x"0757",	
												x"073b",	x"071c",	x"0731",	x"0738",	
												x"072e",	x"0721",	x"0737",	x"0726",	
												x"0746",	x"0739",	x"070d",	x"0743",	
												x"0740",	x"0738",	x"0767",	x"0754",	
												x"0759",	x"0759",	x"075e",	x"075b",	
												x"0755",	x"0741",	x"0750",	x"073d",	
												x"0754",	x"0744",	x"06f9",	x"074b",	
												x"302e",	x"2005",	x"06f4",	x"06da",	
												x"06fe",	x"06e1",	x"06ff",	x"06fd",	
												x"071c",	x"06fe",	x"071d",	x"0719",	
												x"0730",	x"0706",	x"071f",	x"0710",	
												x"06f4",	x"0732",	x"0718",	x"0703",	
												x"0718",	x"0728",	x"0737",	x"071a",	
												x"074c",	x"0729",	x"0730",	x"0726",	
												x"0730",	x"0726",	x"072d",	x"071b",	
												x"06f2",	x"06f6",	x"071c",	x"06fd",	
												x"0734",	x"0733",	x"074e",	x"0743",	
												x"0757",	x"075e",	x"0747",	x"0741",	
												x"0751",	x"0747",	x"073d",	x"073d",	
												x"074a",	x"073d",	x"073e",	x"073c",	
												x"0756",	x"073a",	x"0768",	x"073e",	
												x"076a",	x"072f",	x"0752",	x"073c",	
												x"0759",	x"073c",	x"0763",	x"073a",	
												x"070f",	x"073e",	x"0004",	x"000a",	
												x"3cee",	x"a298",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"2006",	
												x"0713",	x"06e7",	x"0711",	x"0717",	
												x"0747",	x"071d",	x"0747",	x"071a",	
												x"0733",	x"0739",	x"0743",	x"0748",	
												x"074d",	x"074b",	x"0737",	x"0764",	
												x"0745",	x"0746",	x"0763",	x"075b",	
												x"074b",	x"0769",	x"076c",	x"0765",	
												x"076f",	x"074e",	x"076d",	x"0763",	
												x"0779",	x"0786",	x"072a",	x"074c",	
												x"0760",	x"075b",	x"075f",	x"075c",	
												x"0778",	x"0768",	x"077f",	x"0799",	
												x"0777",	x"0770",	x"077d",	x"0780",	
												x"0792",	x"0783",	x"0772",	x"079f",	
												x"079b",	x"0783",	x"0787",	x"078e",	
												x"0798",	x"0784",	x"07c5",	x"079c",	
												x"07b7",	x"07a2",	x"07bd",	x"07a7",	
												x"07b4",	x"07a0",	x"072b",	x"0797",	
												x"502e",	x"2006",	x"0753",	x"073e",	
												x"074f",	x"0731",	x"0763",	x"071e",	
												x"0783",	x"0761",	x"0783",	x"0785",	
												x"0787",	x"0777",	x"0791",	x"076d",	
												x"079a",	x"0764",	x"079b",	x"0799",	
												x"07ae",	x"0788",	x"07a2",	x"078b",	
												x"07a1",	x"07a7",	x"07b3",	x"0797",	
												x"07ab",	x"079e",	x"07a7",	x"07ae",	
												x"077c",	x"0776",	x"07ab",	x"0758",	
												x"07b7",	x"078d",	x"07ba",	x"078e",	
												x"07ea",	x"0789",	x"07da",	x"0790",	
												x"07cc",	x"07a2",	x"07d8",	x"0791",	
												x"0794",	x"0796",	x"07c0",	x"077d",	
												x"07c4",	x"079a",	x"07e0",	x"07a4",	
												x"080a",	x"07a9",	x"07e1",	x"07a4",	
												x"07dd",	x"07a5",	x"07c0",	x"07ae",	
												x"074a",	x"078a",	x"602e",	x"2006",	
												x"0771",	x"073c",	x"078a",	x"071b",	
												x"0785",	x"0780",	x"0798",	x"0772",	
												x"0796",	x"0757",	x"079d",	x"0759",	
												x"078a",	x"07a5",	x"07ab",	x"076e",	
												x"079a",	x"077a",	x"07d2",	x"0777",	
												x"07ce",	x"07a5",	x"07f4",	x"07c4",	
												x"07ea",	x"07b4",	x"07e7",	x"07c3",	
												x"07d1",	x"07b8",	x"07ab",	x"07cb",	
												x"07e1",	x"0788",	x"07e0",	x"07d8",	
												x"07e9",	x"07c3",	x"07f7",	x"07d6",	
												x"07d0",	x"07be",	x"07ec",	x"07d7",	
												x"07e4",	x"07c4",	x"07f7",	x"07d5",	
												x"080c",	x"07b4",	x"080f",	x"07d6",	
												x"080b",	x"07d6",	x"0808",	x"07ef",	
												x"07fb",	x"080a",	x"080e",	x"07ea",	
												x"080a",	x"07b6",	x"0771",	x"07d3",	
												x"702e",	x"2006",	x"0782",	x"0741",	
												x"07c6",	x"075a",	x"07a9",	x"0789",	
												x"0846",	x"07a3",	x"07e8",	x"07a0",	
												x"07ed",	x"07df",	x"07f2",	x"07ec",	
												x"07e4",	x"07e3",	x"0826",	x"07e3",	
												x"082c",	x"081b",	x"082b",	x"080c",	
												x"0877",	x"082f",	x"084f",	x"0811",	
												x"0854",	x"07f1",	x"0832",	x"07f9",	
												x"0810",	x"0822",	x"0852",	x"080a",	
												x"0859",	x"0831",	x"0869",	x"081d",	
												x"085c",	x"0814",	x"0858",	x"0829",	
												x"0862",	x"082b",	x"086b",	x"0831",	
												x"0856",	x"0858",	x"0861",	x"0853",	
												x"086d",	x"085d",	x"0893",	x"084d",	
												x"08ad",	x"0865",	x"08be",	x"086a",	
												x"0896",	x"0863",	x"0867",	x"085d",	
												x"06d8",	x"0864",	x"0004",	x"000a",	
												x"81e2",	x"d872",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"3007",	
												x"06f2",	x"06c2",	x"070c",	x"06e7",	
												x"06dd",	x"0714",	x"06fe",	x"0709",	
												x"06f5",	x"0701",	x"072c",	x"070f",	
												x"071e",	x"0733",	x"06dc",	x"070e",	
												x"0736",	x"070e",	x"073d",	x"071f",	
												x"0743",	x"073e",	x"0756",	x"0745",	
												x"074b",	x"075c",	x"071c",	x"0732",	
												x"070e",	x"0723",	x"0702",	x"0733",	
												x"072a",	x"072a",	x"073f",	x"0732",	
												x"0729",	x"071e",	x"075d",	x"0718",	
												x"072f",	x"073f",	x"0761",	x"073b",	
												x"072f",	x"076a",	x"0702",	x"0730",	
												x"0713",	x"0733",	x"0714",	x"0723",	
												x"0741",	x"0729",	x"0743",	x"074e",	
												x"073f",	x"073f",	x"0757",	x"074a",	
												x"0730",	x"0742",	x"06f3",	x"0717",	
												x"102e",	x"3007",	x"06d3",	x"06d6",	
												x"06e8",	x"06fc",	x"06d9",	x"06d9",	
												x"06ec",	x"06d3",	x"06e7",	x"06e9",	
												x"0703",	x"0704",	x"06f6",	x"0712",	
												x"06f9",	x"0703",	x"071a",	x"070c",	
												x"0715",	x"072a",	x"0709",	x"072e",	
												x"0706",	x"0758",	x"0707",	x"0718",	
												x"0732",	x"06f9",	x"072f",	x"0720",	
												x"070b",	x"073b",	x"0702",	x"072a",	
												x"0700",	x"0706",	x"070a",	x"0700",	
												x"0735",	x"0738",	x"0722",	x"072c",	
												x"073f",	x"0728",	x"0747",	x"0733",	
												x"06f1",	x"0726",	x"0716",	x"0720",	
												x"0726",	x"070f",	x"0727",	x"0742",	
												x"0745",	x"0737",	x"0736",	x"073d",	
												x"0740",	x"072b",	x"0741",	x"073f",	
												x"06d5",	x"0738",	x"202e",	x"3007",	
												x"06ec",	x"06fb",	x"06f1",	x"0700",	
												x"06f1",	x"070b",	x"06e4",	x"070a",	
												x"06dd",	x"071d",	x"071c",	x"06f7",	
												x"0716",	x"073e",	x"06cb",	x"0716",	
												x"0702",	x"06fb",	x"0706",	x"0721",	
												x"0708",	x"0719",	x"0709",	x"0708",	
												x"0715",	x"0719",	x"071e",	x"071d",	
												x"0714",	x"0706",	x"06d9",	x"06f7",	
												x"0704",	x"0705",	x"0709",	x"06f4",	
												x"070e",	x"070f",	x"070e",	x"070d",	
												x"071a",	x"0700",	x"0725",	x"071b",	
												x"072a",	x"0722",	x"06f6",	x"070c",	
												x"06dd",	x"0700",	x"0721",	x"06f2",	
												x"0702",	x"0705",	x"071a",	x"0716",	
												x"0711",	x"072b",	x"072b",	x"0713",	
												x"0736",	x"0715",	x"06cd",	x"071f",	
												x"302e",	x"3007",	x"06cf",	x"06aa",	
												x"06dc",	x"06c5",	x"06d8",	x"06d0",	
												x"06ef",	x"06f5",	x"06e3",	x"06c3",	
												x"06d3",	x"06d5",	x"06d4",	x"06d3",	
												x"06cb",	x"06d8",	x"06fb",	x"06e2",	
												x"06f3",	x"06f1",	x"0703",	x"06e7",	
												x"0703",	x"0710",	x"0723",	x"06f9",	
												x"070c",	x"070a",	x"0710",	x"0710",	
												x"06e4",	x"070d",	x"06fb",	x"06de",	
												x"06f6",	x"06f0",	x"0707",	x"06e5",	
												x"070c",	x"0718",	x"0724",	x"070e",	
												x"0725",	x"072d",	x"0716",	x"0715",	
												x"0708",	x"0709",	x"0712",	x"070d",	
												x"06fa",	x"0727",	x"0709",	x"06e1",	
												x"0746",	x"0710",	x"0739",	x"070d",	
												x"0746",	x"0728",	x"071d",	x"06fd",	
												x"06e7",	x"0707",	x"0004",	x"000a",	
												x"2704",	x"ccf7",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"3008",	
												x"06e1",	x"06bb",	x"06cc",	x"06d4",	
												x"06ef",	x"06ea",	x"06d4",	x"0705",	
												x"06ee",	x"06ee",	x"0707",	x"06e5",	
												x"0711",	x"070f",	x"06eb",	x"070b",	
												x"0721",	x"0720",	x"0702",	x"072b",	
												x"072e",	x"0712",	x"073a",	x"0736",	
												x"0732",	x"0735",	x"0740",	x"072c",	
												x"071c",	x"0747",	x"0706",	x"0707",	
												x"072d",	x"0716",	x"0721",	x"0722",	
												x"073d",	x"071e",	x"0747",	x"0732",	
												x"075c",	x"072c",	x"0757",	x"0748",	
												x"0761",	x"073d",	x"0708",	x"0743",	
												x"0745",	x"0742",	x"0751",	x"073f",	
												x"075b",	x"0758",	x"0763",	x"076c",	
												x"0769",	x"074f",	x"077f",	x"0769",	
												x"0766",	x"0756",	x"0710",	x"075b",	
												x"502e",	x"3008",	x"0703",	x"06ec",	
												x"072f",	x"06f2",	x"0730",	x"06fb",	
												x"0738",	x"0728",	x"0738",	x"070a",	
												x"070f",	x"071c",	x"074e",	x"072f",	
												x"0753",	x"0756",	x"0757",	x"0729",	
												x"075e",	x"0768",	x"0753",	x"077c",	
												x"076b",	x"075d",	x"0777",	x"0755",	
												x"0773",	x"0766",	x"0763",	x"0764",	
												x"074b",	x"0748",	x"0751",	x"071a",	
												x"075b",	x"072a",	x"076a",	x"074b",	
												x"07ae",	x"0768",	x"0792",	x"078a",	
												x"079b",	x"0768",	x"0799",	x"0778",	
												x"0766",	x"077a",	x"0796",	x"0748",	
												x"0777",	x"076f",	x"0793",	x"075f",	
												x"079d",	x"0772",	x"07a3",	x"076b",	
												x"07a4",	x"0783",	x"078b",	x"0768",	
												x"072b",	x"0760",	x"602e",	x"3008",	
												x"0736",	x"0718",	x"072f",	x"071d",	
												x"072c",	x"074c",	x"071c",	x"070d",	
												x"0751",	x"0730",	x"0746",	x"0766",	
												x"0768",	x"0751",	x"0762",	x"0754",	
												x"0791",	x"0765",	x"0791",	x"0775",	
												x"078d",	x"0783",	x"0797",	x"0786",	
												x"0791",	x"0772",	x"0794",	x"077f",	
												x"0792",	x"0783",	x"0754",	x"0780",	
												x"0783",	x"0765",	x"0796",	x"079c",	
												x"07ad",	x"078d",	x"07d6",	x"0783",	
												x"07c6",	x"07af",	x"07c3",	x"07b2",	
												x"07b4",	x"0788",	x"07a6",	x"079a",	
												x"07c5",	x"07a3",	x"0796",	x"07ac",	
												x"07c7",	x"076c",	x"07f7",	x"07aa",	
												x"07e9",	x"07c8",	x"07e8",	x"07ce",	
												x"07cf",	x"07bf",	x"0755",	x"07a8",	
												x"702e",	x"3008",	x"078c",	x"0735",	
												x"0785",	x"0774",	x"0759",	x"0756",	
												x"07aa",	x"0748",	x"0780",	x"078e",	
												x"078e",	x"0779",	x"07a7",	x"077e",	
												x"07ac",	x"07a5",	x"07e1",	x"07b1",	
												x"07e9",	x"07c5",	x"07f4",	x"07bb",	
												x"07f6",	x"07bb",	x"0813",	x"07c3",	
												x"07fc",	x"080c",	x"07f7",	x"07f6",	
												x"07dd",	x"07fd",	x"07fd",	x"07dd",	
												x"0806",	x"07fd",	x"080a",	x"07ea",	
												x"0832",	x"07e3",	x"0812",	x"07fb",	
												x"083c",	x"083e",	x"0805",	x"081b",	
												x"0817",	x"0818",	x"080b",	x"0831",	
												x"082a",	x"07ce",	x"082e",	x"07f1",	
												x"0880",	x"082c",	x"0878",	x"082f",	
												x"0877",	x"084a",	x"0832",	x"0840",	
												x"06cc",	x"0816",	x"0004",	x"000a",	
												x"60dc",	x"fd30",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"0009",	
												x"06d3",	x"06d9",	x"06fa",	x"06f4",	
												x"06c7",	x"06fd",	x"06e3",	x"06d1",	
												x"06e6",	x"06cf",	x"069a",	x"06d3",	
												x"0691",	x"06b3",	x"066e",	x"0684",	
												x"069f",	x"0694",	x"06c5",	x"06b9",	
												x"06bf",	x"06c4",	x"06c5",	x"06cf",	
												x"06de",	x"06cf",	x"0715",	x"0708",	
												x"0713",	x"06f9",	x"06ad",	x"06e7",	
												x"06d0",	x"06c9",	x"06ca",	x"06c5",	
												x"06df",	x"06d1",	x"06e8",	x"06f6",	
												x"06f2",	x"06c6",	x"0708",	x"06f9",	
												x"0710",	x"070f",	x"06a7",	x"06e9",	
												x"06d8",	x"06cb",	x"06ea",	x"06c1",	
												x"06f7",	x"06c5",	x"06e7",	x"06f4",	
												x"0701",	x"06d9",	x"0742",	x"06f9",	
												x"072d",	x"0708",	x"06bb",	x"06f5",	
												x"102f",	x"0009",	x"06c4",	x"06e3",	
												x"06ed",	x"06b1",	x"06a8",	x"06ba",	
												x"06ce",	x"069e",	x"069f",	x"06a4",	
												x"06a1",	x"06c6",	x"066f",	x"0699",	
												x"0667",	x"06a4",	x"06a3",	x"0655",	
												x"06c5",	x"06a9",	x"06be",	x"0690",	
												x"06cf",	x"06cb",	x"06e2",	x"06d7",	
												x"06fb",	x"06e4",	x"06f5",	x"06ec",	
												x"06ad",	x"06e1",	x"06a5",	x"06bf",	
												x"06d4",	x"06fc",	x"06d2",	x"06c2",	
												x"06e1",	x"06ec",	x"06d4",	x"06ef",	
												x"06c1",	x"06e8",	x"06cb",	x"06be",	
												x"06b9",	x"06b8",	x"06d4",	x"06d7",	
												x"06c6",	x"06e9",	x"06d9",	x"06db",	
												x"06e4",	x"06df",	x"0708",	x"06dd",	
												x"0720",	x"0700",	x"0713",	x"06f7",	
												x"069e",	x"070d",	x"202f",	x"0009",	
												x"06ad",	x"069f",	x"068a",	x"069c",	
												x"06b8",	x"0680",	x"0696",	x"06a4",	
												x"0695",	x"0671",	x"0674",	x"06a5",	
												x"0677",	x"0699",	x"0622",	x"0683",	
												x"068c",	x"0662",	x"06bd",	x"06ab",	
												x"06c2",	x"06a9",	x"06c9",	x"06cb",	
												x"06dd",	x"06ca",	x"06e5",	x"06ea",	
												x"06db",	x"06d5",	x"06c6",	x"06d1",	
												x"06b0",	x"06b4",	x"06d1",	x"06b8",	
												x"06cb",	x"06d2",	x"06d8",	x"06e7",	
												x"06dd",	x"06cb",	x"06d8",	x"06d9",	
												x"06f0",	x"06c7",	x"06b7",	x"06ee",	
												x"06d7",	x"06f3",	x"06d4",	x"06b8",	
												x"06cc",	x"06c2",	x"06c9",	x"06ce",	
												x"06f8",	x"06c1",	x"06fe",	x"06e6",	
												x"0702",	x"06e4",	x"069c",	x"06dd",	
												x"302f",	x"0009",	x"06b6",	x"065e",	
												x"0698",	x"06a3",	x"06a0",	x"068a",	
												x"069a",	x"0673",	x"06c7",	x"067e",	
												x"06a9",	x"06a1",	x"0697",	x"06a0",	
												x"0682",	x"0696",	x"06a9",	x"0656",	
												x"06b2",	x"068a",	x"06ce",	x"06a9",	
												x"06e8",	x"0695",	x"06e8",	x"06c6",	
												x"06cd",	x"06c6",	x"06d7",	x"06d1",	
												x"0697",	x"06c7",	x"06c4",	x"06a4",	
												x"06ce",	x"06af",	x"06d0",	x"06bb",	
												x"06e3",	x"06d0",	x"06e9",	x"06ce",	
												x"06e2",	x"06ec",	x"0714",	x"06d2",	
												x"06a9",	x"06cf",	x"06f5",	x"06cc",	
												x"06ea",	x"06d5",	x"06f3",	x"06ae",	
												x"0711",	x"06d8",	x"0734",	x"06d3",	
												x"071e",	x"06e5",	x"0728",	x"06fc",	
												x"06b0",	x"06e8",	x"0004",	x"000a",	
												x"05fd",	x"e6e1",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"000a",	
												x"06c4",	x"069e",	x"06cc",	x"06a2",	
												x"06e1",	x"068a",	x"06f0",	x"06b1",	
												x"06c2",	x"06ad",	x"06ce",	x"069f",	
												x"06b8",	x"0693",	x"0688",	x"06a5",	
												x"06f6",	x"0676",	x"06ef",	x"06be",	
												x"0728",	x"06bd",	x"0731",	x"06d8",	
												x"0709",	x"06e1",	x"070d",	x"06f8",	
												x"0714",	x"0709",	x"06ed",	x"06f7",	
												x"0723",	x"06f7",	x"071d",	x"0706",	
												x"071f",	x"06f7",	x"0734",	x"0703",	
												x"0732",	x"0710",	x"0730",	x"0722",	
												x"0742",	x"0721",	x"070f",	x"0700",	
												x"0744",	x"0705",	x"073b",	x"071a",	
												x"0737",	x"06dc",	x"075d",	x"072c",	
												x"0763",	x"071a",	x"075e",	x"071f",	
												x"0747",	x"0713",	x"06e2",	x"0711",	
												x"502f",	x"000a",	x"0703",	x"06dd",	
												x"0717",	x"06df",	x"06f8",	x"06e2",	
												x"0707",	x"06dd",	x"06fd",	x"06e3",	
												x"0710",	x"06e7",	x"070f",	x"06b7",	
												x"06de",	x"06ce",	x"0737",	x"06ce",	
												x"0724",	x"06d8",	x"073c",	x"06c0",	
												x"0745",	x"070d",	x"0748",	x"071a",	
												x"074c",	x"0742",	x"0740",	x"0704",	
												x"0734",	x"0718",	x"0750",	x"06ef",	
												x"0763",	x"071e",	x"074e",	x"06eb",	
												x"0759",	x"0721",	x"0773",	x"071f",	
												x"076b",	x"073d",	x"0756",	x"073f",	
												x"0745",	x"0710",	x"0781",	x"0712",	
												x"0776",	x"072c",	x"0778",	x"071f",	
												x"0787",	x"071f",	x"0791",	x"072f",	
												x"079e",	x"0752",	x"0783",	x"074b",	
												x"06d5",	x"073c",	x"602f",	x"000a",	
												x"0709",	x"06b7",	x"06fd",	x"06df",	
												x"073f",	x"06e4",	x"071c",	x"06fa",	
												x"0705",	x"06f3",	x"0704",	x"06d7",	
												x"0703",	x"06c7",	x"06fc",	x"06f3",	
												x"0723",	x"06c3",	x"074a",	x"06f4",	
												x"075d",	x"0728",	x"0773",	x"0720",	
												x"077c",	x"0737",	x"0782",	x"0740",	
												x"077d",	x"074e",	x"0756",	x"0740",	
												x"079a",	x"072e",	x"0791",	x"0744",	
												x"079d",	x"0745",	x"07a0",	x"0758",	
												x"0780",	x"074e",	x"0794",	x"0767",	
												x"07a0",	x"074a",	x"0765",	x"077c",	
												x"0790",	x"0754",	x"07c0",	x"0751",	
												x"07b1",	x"0777",	x"0813",	x"0760",	
												x"07ea",	x"0769",	x"07c6",	x"07a6",	
												x"07cf",	x"0785",	x"0739",	x"0789",	
												x"702f",	x"000a",	x"073a",	x"06f8",	
												x"0757",	x"0707",	x"0735",	x"06f9",	
												x"0767",	x"0707",	x"074a",	x"0713",	
												x"077a",	x"06fb",	x"074a",	x"0721",	
												x"0721",	x"0710",	x"0785",	x"06e9",	
												x"07a7",	x"0739",	x"07dc",	x"0759",	
												x"07e4",	x"074f",	x"07d4",	x"0771",	
												x"07cc",	x"0785",	x"07ec",	x"0796",	
												x"0782",	x"078f",	x"07e0",	x"0781",	
												x"07dd",	x"07a2",	x"07ed",	x"079a",	
												x"07f1",	x"078f",	x"07fb",	x"0779",	
												x"07e9",	x"07d3",	x"080c",	x"0793",	
												x"07b1",	x"07bd",	x"07ed",	x"0793",	
												x"0805",	x"07bf",	x"081e",	x"07c0",	
												x"0829",	x"07be",	x"082a",	x"07d5",	
												x"083a",	x"07eb",	x"081a",	x"07ff",	
												x"0683",	x"07d5",	x"0004",	x"000a",	
												x"4e38",	x"1612",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"100b",	
												x"069d",	x"067e",	x"06bd",	x"0693",	
												x"0694",	x"06ab",	x"0663",	x"0677",	
												x"066b",	x"0645",	x"0670",	x"064c",	
												x"065f",	x"063b",	x"064e",	x"0637",	
												x"0675",	x"0669",	x"0673",	x"069c",	
												x"0691",	x"067b",	x"0685",	x"06ab",	
												x"06a9",	x"068e",	x"06a6",	x"06c6",	
												x"069c",	x"069e",	x"066f",	x"06ba",	
												x"068d",	x"0681",	x"06b9",	x"06a4",	
												x"0685",	x"067d",	x"0699",	x"068f",	
												x"06a4",	x"068f",	x"06a1",	x"0699",	
												x"0687",	x"06a7",	x"066c",	x"06a2",	
												x"06a4",	x"0684",	x"069c",	x"06a1",	
												x"0684",	x"0689",	x"06a9",	x"0667",	
												x"06b3",	x"06b7",	x"06ba",	x"069a",	
												x"06b3",	x"0694",	x"0670",	x"0699",	
												x"102f",	x"100b",	x"067a",	x"0655",	
												x"0688",	x"0661",	x"064d",	x"0686",	
												x"0652",	x"0658",	x"0636",	x"061e",	
												x"0633",	x"0621",	x"0624",	x"062b",	
												x"0631",	x"0675",	x"064e",	x"0628",	
												x"067c",	x"0640",	x"06bc",	x"0661",	
												x"0694",	x"0688",	x"0698",	x"0687",	
												x"0687",	x"069f",	x"068d",	x"068b",	
												x"0649",	x"069a",	x"0674",	x"0658",	
												x"0668",	x"0666",	x"068f",	x"0683",	
												x"067e",	x"06a3",	x"06a2",	x"066e",	
												x"0693",	x"06a9",	x"06a5",	x"06a0",	
												x"0657",	x"0694",	x"0687",	x"066b",	
												x"06a2",	x"069b",	x"06b4",	x"0697",	
												x"06b7",	x"06ac",	x"06c8",	x"06af",	
												x"06c3",	x"06b7",	x"06a9",	x"06b7",	
												x"0657",	x"06a2",	x"202f",	x"100b",	
												x"0665",	x"065f",	x"0680",	x"066b",	
												x"0653",	x"0655",	x"0652",	x"0640",	
												x"0625",	x"0647",	x"0645",	x"0638",	
												x"0629",	x"063f",	x"061a",	x"0642",	
												x"0632",	x"063e",	x"0659",	x"064e",	
												x"0662",	x"066b",	x"067d",	x"0686",	
												x"0688",	x"069c",	x"0698",	x"068a",	
												x"0681",	x"067c",	x"0658",	x"067b",	
												x"066c",	x"0652",	x"068b",	x"0676",	
												x"067a",	x"068b",	x"0679",	x"0675",	
												x"0682",	x"0676",	x"068b",	x"0681",	
												x"0686",	x"0667",	x"0669",	x"0687",	
												x"0669",	x"068c",	x"0684",	x"0680",	
												x"0685",	x"0673",	x"068c",	x"067e",	
												x"0690",	x"066c",	x"069c",	x"068c",	
												x"069b",	x"0687",	x"066a",	x"0675",	
												x"302f",	x"100b",	x"0663",	x"065a",	
												x"0662",	x"0636",	x"0663",	x"0632",	
												x"0641",	x"0631",	x"063f",	x"062a",	
												x"063e",	x"0620",	x"0644",	x"0629",	
												x"0639",	x"064a",	x"0622",	x"0628",	
												x"0663",	x"0640",	x"0676",	x"063d",	
												x"069d",	x"0660",	x"068b",	x"0672",	
												x"06a2",	x"0673",	x"068f",	x"0687",	
												x"0669",	x"065a",	x"0678",	x"065c",	
												x"067d",	x"066e",	x"0678",	x"0662",	
												x"0684",	x"0680",	x"0696",	x"0681",	
												x"06a4",	x"0681",	x"068b",	x"0685",	
												x"0693",	x"0678",	x"0694",	x"067d",	
												x"06a2",	x"0672",	x"0693",	x"0668",	
												x"0694",	x"067c",	x"06b0",	x"0679",	
												x"06c0",	x"0683",	x"06ab",	x"0682",	
												x"0667",	x"068b",	x"0004",	x"000a",	
												x"de00",	x"fe3b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"100c",	
												x"067b",	x"0630",	x"0690",	x"065e",	
												x"066f",	x"0659",	x"0672",	x"0670",	
												x"0663",	x"0654",	x"066e",	x"0656",	
												x"0659",	x"063e",	x"066e",	x"065c",	
												x"0679",	x"0635",	x"068b",	x"063f",	
												x"06b1",	x"0678",	x"06be",	x"0691",	
												x"06c0",	x"06a1",	x"06cf",	x"06a6",	
												x"06a7",	x"06a5",	x"06ae",	x"0680",	
												x"06d3",	x"0697",	x"06d2",	x"06be",	
												x"06d0",	x"06b6",	x"06d5",	x"06d0",	
												x"06ca",	x"06cc",	x"06df",	x"06bb",	
												x"06be",	x"06ce",	x"06b9",	x"06b4",	
												x"06d5",	x"06c0",	x"06d3",	x"06ac",	
												x"06df",	x"06b8",	x"06eb",	x"06c4",	
												x"0700",	x"06c6",	x"06f0",	x"06e4",	
												x"0701",	x"06bf",	x"0698",	x"06dc",	
												x"502f",	x"100c",	x"0688",	x"0685",	
												x"0688",	x"0678",	x"0697",	x"067a",	
												x"06a5",	x"0685",	x"06a6",	x"0685",	
												x"06c0",	x"0683",	x"06b0",	x"06b1",	
												x"0694",	x"0682",	x"06e1",	x"068d",	
												x"06cb",	x"06aa",	x"06d1",	x"0684",	
												x"06fb",	x"06cc",	x"0707",	x"06b4",	
												x"06ea",	x"06c5",	x"06f7",	x"06bb",	
												x"06c7",	x"06cd",	x"06d3",	x"069c",	
												x"0702",	x"06b9",	x"0713",	x"06bc",	
												x"0713",	x"06da",	x"070c",	x"06d3",	
												x"0701",	x"06e6",	x"0705",	x"06e6",	
												x"06f6",	x"06d6",	x"06f2",	x"06d1",	
												x"070f",	x"06c0",	x"072d",	x"06db",	
												x"0731",	x"06dc",	x"072f",	x"06ed",	
												x"072e",	x"06fe",	x"0715",	x"06f5",	
												x"06ae",	x"06ea",	x"602f",	x"100c",	
												x"06c3",	x"068d",	x"06d5",	x"0677",	
												x"06a9",	x"0682",	x"06a5",	x"0670",	
												x"06cd",	x"067a",	x"06a9",	x"066a",	
												x"06a6",	x"0671",	x"06a9",	x"0680",	
												x"06b7",	x"0693",	x"06c4",	x"069b",	
												x"070f",	x"0699",	x"0722",	x"06e9",	
												x"071f",	x"06f2",	x"0710",	x"06fe",	
												x"06ff",	x"06d9",	x"06e2",	x"06d3",	
												x"072d",	x"06c5",	x"0717",	x"0726",	
												x"072c",	x"06ff",	x"0736",	x"0708",	
												x"073b",	x"06f5",	x"0742",	x"0708",	
												x"0741",	x"071c",	x"072e",	x"06fe",	
												x"072f",	x"0700",	x"0724",	x"0709",	
												x"074c",	x"06fb",	x"073a",	x"070f",	
												x"0762",	x"0710",	x"074e",	x"072a",	
												x"0737",	x"072b",	x"06f8",	x"071d",	
												x"702f",	x"100c",	x"06d4",	x"0686",	
												x"06d0",	x"069b",	x"06f1",	x"06b5",	
												x"06d9",	x"06c5",	x"06e3",	x"066f",	
												x"06f2",	x"06c5",	x"06e3",	x"06b0",	
												x"06c3",	x"06ce",	x"072d",	x"069e",	
												x"0726",	x"0702",	x"0744",	x"0718",	
												x"075f",	x"0728",	x"0762",	x"071a",	
												x"077e",	x"0759",	x"0735",	x"0712",	
												x"0728",	x"071b",	x"0773",	x"06ee",	
												x"0766",	x"0726",	x"077b",	x"0725",	
												x"0795",	x"076d",	x"07a2",	x"0750",	
												x"0791",	x"074f",	x"078e",	x"0747",	
												x"075a",	x"075a",	x"0798",	x"074f",	
												x"07ad",	x"076a",	x"0798",	x"0753",	
												x"07ca",	x"0773",	x"07c3",	x"0787",	
												x"07b7",	x"079b",	x"07ae",	x"079f",	
												x"0703",	x"0771",	x"0004",	x"000a",	
												x"1d1a",	x"2bff",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"200d",	
												x"072c",	x"0716",	x"0729",	x"0760",	
												x"070a",	x"0720",	x"0730",	x"0721",	
												x"0728",	x"0725",	x"0713",	x"06f5",	
												x"0738",	x"0709",	x"071e",	x"074d",	
												x"0771",	x"0752",	x"0773",	x"0768",	
												x"075d",	x"0778",	x"0762",	x"0777",	
												x"0766",	x"0764",	x"0799",	x"0773",	
												x"0757",	x"077d",	x"0716",	x"072d",	
												x"0751",	x"0739",	x"0746",	x"0786",	
												x"0745",	x"0761",	x"0756",	x"0767",	
												x"0759",	x"0760",	x"075c",	x"0764",	
												x"0771",	x"0768",	x"0748",	x"076d",	
												x"076c",	x"076c",	x"07a4",	x"0778",	
												x"0787",	x"0781",	x"0759",	x"076a",	
												x"076c",	x"0766",	x"0779",	x"0761",	
												x"0779",	x"0764",	x"06ec",	x"075f",	
												x"102f",	x"200d",	x"0719",	x"070a",	
												x"0738",	x"0710",	x"0702",	x"0741",	
												x"06fd",	x"071b",	x"06f4",	x"06db",	
												x"0713",	x"0715",	x"071b",	x"0735",	
												x"06e4",	x"0729",	x"073a",	x"0711",	
												x"074f",	x"0731",	x"0760",	x"0772",	
												x"075e",	x"076c",	x"0754",	x"074b",	
												x"0764",	x"0760",	x"075d",	x"076a",	
												x"070b",	x"0759",	x"071f",	x"070a",	
												x"073f",	x"072f",	x"075b",	x"0745",	
												x"0768",	x"075c",	x"0730",	x"075a",	
												x"076e",	x"0750",	x"0758",	x"074a",	
												x"0749",	x"0767",	x"075a",	x"0760",	
												x"075f",	x"075b",	x"078a",	x"075e",	
												x"0763",	x"0776",	x"0766",	x"075d",	
												x"0770",	x"0755",	x"0764",	x"0752",	
												x"06fe",	x"075a",	x"202f",	x"200d",	
												x"0714",	x"0720",	x"06fa",	x"0713",	
												x"0705",	x"0706",	x"06fa",	x"071e",	
												x"06f9",	x"06f0",	x"06fa",	x"071f",	
												x"0744",	x"0716",	x"06e8",	x"0734",	
												x"0721",	x"070c",	x"0757",	x"073c",	
												x"0748",	x"0746",	x"0754",	x"074d",	
												x"073d",	x"073d",	x"0750",	x"0746",	
												x"074e",	x"0746",	x"0712",	x"0736",	
												x"073e",	x"0706",	x"074a",	x"0762",	
												x"0734",	x"073a",	x"0731",	x"0739",	
												x"073a",	x"073e",	x"0754",	x"0737",	
												x"074d",	x"0750",	x"0748",	x"074e",	
												x"075c",	x"0757",	x"0756",	x"0746",	
												x"075a",	x"073d",	x"074c",	x"0754",	
												x"0754",	x"0726",	x"074a",	x"0749",	
												x"075f",	x"073c",	x"06cc",	x"0755",	
												x"302f",	x"200d",	x"070c",	x"06b7",	
												x"071d",	x"06ff",	x"070b",	x"06fb",	
												x"06ef",	x"06fb",	x"06f1",	x"06d0",	
												x"071d",	x"06d3",	x"070f",	x"06e3",	
												x"0708",	x"0707",	x"072f",	x"06f7",	
												x"0760",	x"0730",	x"0754",	x"0744",	
												x"0748",	x"0746",	x"0749",	x"0741",	
												x"0744",	x"0750",	x"0743",	x"072f",	
												x"0713",	x"0718",	x"0755",	x"0722",	
												x"073e",	x"074c",	x"0744",	x"0740",	
												x"0763",	x"0746",	x"077f",	x"074c",	
												x"0795",	x"075b",	x"076d",	x"0750",	
												x"076a",	x"075a",	x"0777",	x"074a",	
												x"076b",	x"0748",	x"077e",	x"074f",	
												x"0777",	x"073c",	x"077d",	x"0748",	
												x"0784",	x"0769",	x"0783",	x"0747",	
												x"070d",	x"074f",	x"0004",	x"000a",	
												x"40dd",	x"a372",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"200e",	
												x"0749",	x"0707",	x"0729",	x"070d",	
												x"0710",	x"06f2",	x"0715",	x"06e4",	
												x"072a",	x"06f7",	x"072d",	x"072c",	
												x"0773",	x"0725",	x"074f",	x"0739",	
												x"0769",	x"075b",	x"0776",	x"0779",	
												x"0761",	x"0760",	x"076c",	x"076d",	
												x"0786",	x"0765",	x"0775",	x"076c",	
												x"0771",	x"0775",	x"0773",	x"075f",	
												x"078b",	x"0759",	x"0780",	x"0783",	
												x"079a",	x"0771",	x"07b4",	x"0775",	
												x"07b6",	x"075d",	x"07ae",	x"0793",	
												x"07bb",	x"078d",	x"0792",	x"07ae",	
												x"07c1",	x"078f",	x"07b4",	x"07b2",	
												x"07c7",	x"07a0",	x"07af",	x"07a1",	
												x"07c2",	x"0790",	x"07d8",	x"07b2",	
												x"07d7",	x"07a8",	x"0769",	x"0797",	
												x"502f",	x"200e",	x"077f",	x"0739",	
												x"0794",	x"0771",	x"077d",	x"0740",	
												x"0775",	x"0756",	x"0758",	x"0719",	
												x"079a",	x"072c",	x"078b",	x"0777",	
												x"0788",	x"073c",	x"07a1",	x"0795",	
												x"07c2",	x"076b",	x"07d6",	x"0791",	
												x"07c9",	x"07a2",	x"07b4",	x"079c",	
												x"07a2",	x"079a",	x"07d7",	x"07a3",	
												x"0798",	x"078a",	x"07cf",	x"077b",	
												x"07d1",	x"07c1",	x"07dc",	x"0796",	
												x"07ea",	x"07ab",	x"07e2",	x"07a4",	
												x"07f3",	x"07a7",	x"07fe",	x"07a7",	
												x"07c7",	x"07aa",	x"080b",	x"0799",	
												x"07d2",	x"07a9",	x"07e9",	x"07a6",	
												x"07f9",	x"07a8",	x"0814",	x"07a6",	
												x"080e",	x"07c6",	x"0801",	x"07ba",	
												x"075d",	x"07a4",	x"602f",	x"200e",	
												x"0786",	x"0738",	x"0782",	x"076b",	
												x"077e",	x"0768",	x"079b",	x"074e",	
												x"078c",	x"0764",	x"077d",	x"0765",	
												x"078b",	x"0760",	x"0797",	x"0769",	
												x"07fe",	x"075d",	x"0802",	x"079c",	
												x"0813",	x"07aa",	x"0819",	x"07cf",	
												x"07ec",	x"07aa",	x"07d6",	x"07b4",	
												x"07ce",	x"07bd",	x"07d2",	x"07c3",	
												x"07e4",	x"07b2",	x"080c",	x"07c0",	
												x"0821",	x"07b5",	x"080c",	x"07d3",	
												x"0833",	x"07c4",	x"083b",	x"0812",	
												x"082b",	x"07e6",	x"07fc",	x"07bd",	
												x"082a",	x"07d8",	x"081e",	x"07d0",	
												x"085c",	x"07ce",	x"082b",	x"07e7",	
												x"084f",	x"07e3",	x"0834",	x"0811",	
												x"0841",	x"07e7",	x"07b3",	x"07d8",	
												x"702f",	x"200e",	x"07d8",	x"076a",	
												x"0789",	x"0770",	x"07c4",	x"076e",	
												x"07e9",	x"077d",	x"07bd",	x"0786",	
												x"07d4",	x"0768",	x"07ec",	x"0775",	
												x"07fd",	x"07aa",	x"0845",	x"07f1",	
												x"084b",	x"0804",	x"0862",	x"0803",	
												x"0853",	x"0811",	x"0850",	x"0807",	
												x"0876",	x"0801",	x"083f",	x"0839",	
												x"0847",	x"0801",	x"0849",	x"0812",	
												x"082c",	x"080e",	x"0891",	x"0809",	
												x"0897",	x"082f",	x"088e",	x"0823",	
												x"0885",	x"084b",	x"088c",	x"0860",	
												x"084d",	x"0851",	x"088e",	x"0841",	
												x"0888",	x"085f",	x"08ba",	x"0858",	
												x"0899",	x"0887",	x"08b0",	x"0854",	
												x"08b0",	x"0856",	x"08ad",	x"086a",	
												x"0743",	x"0852",	x"0004",	x"000a",	
												x"8ddf",	x"d841",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"300f",	
												x"06ec",	x"0710",	x"06fb",	x"0705",	
												x"06ea",	x"06ee",	x"06e2",	x"06f4",	
												x"06e6",	x"06f0",	x"06fd",	x"06f3",	
												x"0711",	x"06ed",	x"06fa",	x"0746",	
												x"0739",	x"06fd",	x"0735",	x"073a",	
												x"0746",	x"0752",	x"076d",	x"0759",	
												x"0764",	x"075c",	x"074e",	x"0761",	
												x"0728",	x"0763",	x"06f4",	x"074c",	
												x"072b",	x"0727",	x"0733",	x"0740",	
												x"0721",	x"073c",	x"0734",	x"073a",	
												x"077f",	x"071b",	x"076c",	x"0763",	
												x"074f",	x"0758",	x"0707",	x"073e",	
												x"074c",	x"0748",	x"0749",	x"0756",	
												x"0741",	x"071c",	x"074a",	x"0733",	
												x"073f",	x"072e",	x"0779",	x"0749",	
												x"076a",	x"074f",	x"06d4",	x"0753",	
												x"102f",	x"300f",	x"06e7",	x"06d4",	
												x"06f6",	x"06fe",	x"06c3",	x"06e9",	
												x"06c2",	x"06c4",	x"06c3",	x"06dd",	
												x"06ec",	x"06eb",	x"0703",	x"06e2",	
												x"06f0",	x"06d7",	x"06ff",	x"06f3",	
												x"0741",	x"0722",	x"0740",	x"074b",	
												x"075a",	x"0760",	x"0736",	x"073b",	
												x"072a",	x"0749",	x"0702",	x"0723",	
												x"06e5",	x"070f",	x"06ec",	x"06fa",	
												x"070b",	x"0708",	x"0732",	x"06f8",	
												x"0738",	x"0752",	x"071f",	x"0729",	
												x"071c",	x"0744",	x"074a",	x"0727",	
												x"0716",	x"0735",	x"072e",	x"0751",	
												x"0754",	x"0754",	x"073e",	x"0723",	
												x"0726",	x"071e",	x"072c",	x"071d",	
												x"0744",	x"073b",	x"074a",	x"073f",	
												x"06f2",	x"0761",	x"202f",	x"300f",	
												x"06e4",	x"06d6",	x"06d6",	x"06d8",	
												x"06f2",	x"06d6",	x"06d1",	x"06fe",	
												x"06d7",	x"06ec",	x"06f9",	x"06e0",	
												x"06ac",	x"06f5",	x"06a0",	x"06db",	
												x"06f2",	x"06f9",	x"0718",	x"0731",	
												x"0720",	x"0724",	x"0714",	x"070a",	
												x"0713",	x"071b",	x"070e",	x"0729",	
												x"070a",	x"0701",	x"06cb",	x"0707",	
												x"0711",	x"06ee",	x"070a",	x"0726",	
												x"0702",	x"06f3",	x"070d",	x"070b",	
												x"0725",	x"0709",	x"0739",	x"0718",	
												x"0737",	x"073b",	x"0712",	x"0721",	
												x"0724",	x"0725",	x"072d",	x"0722",	
												x"0736",	x"071f",	x"0732",	x"0724",	
												x"071b",	x"071d",	x"0726",	x"070e",	
												x"073e",	x"0714",	x"06e1",	x"0710",	
												x"302f",	x"300f",	x"06f6",	x"06c9",	
												x"06da",	x"06d2",	x"06c6",	x"06cd",	
												x"06cf",	x"06ac",	x"06d3",	x"06a7",	
												x"06c6",	x"06c6",	x"06e2",	x"06c7",	
												x"06c0",	x"06c3",	x"0701",	x"06d3",	
												x"071a",	x"070c",	x"0717",	x"06f3",	
												x"0726",	x"0719",	x"072d",	x"0702",	
												x"072e",	x"071b",	x"0706",	x"070a",	
												x"06e3",	x"06f9",	x"0720",	x"06d8",	
												x"071b",	x"071c",	x"072b",	x"06f3",	
												x"0725",	x"072b",	x"071e",	x"071b",	
												x"073f",	x"0719",	x"073c",	x"071e",	
												x"0740",	x"0712",	x"0741",	x"0722",	
												x"072a",	x"072e",	x"071d",	x"0700",	
												x"072b",	x"070b",	x"0730",	x"0705",	
												x"0749",	x"0702",	x"073d",	x"0701",	
												x"06f7",	x"070e",	x"0004",	x"000a",	
												x"2a9c",	x"ce0d",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"3010",	
												x"06e6",	x"06d3",	x"06e3",	x"06d0",	
												x"06ee",	x"06de",	x"06fe",	x"06fa",	
												x"0708",	x"06f0",	x"06f9",	x"06ec",	
												x"072a",	x"06f4",	x"0707",	x"071f",	
												x"073d",	x"06ed",	x"0732",	x"0730",	
												x"0732",	x"072c",	x"074d",	x"072c",	
												x"0751",	x"072f",	x"074a",	x"0731",	
												x"0733",	x"0726",	x"0713",	x"0701",	
												x"0754",	x"0711",	x"076d",	x"074b",	
												x"0769",	x"0744",	x"0776",	x"0754",	
												x"0776",	x"074f",	x"0775",	x"075b",	
												x"0788",	x"075d",	x"074f",	x"0759",	
												x"076c",	x"0760",	x"0770",	x"0763",	
												x"075d",	x"075b",	x"078e",	x"0761",	
												x"0788",	x"0755",	x"0795",	x"0765",	
												x"0782",	x"075e",	x"072e",	x"074b",	
												x"502f",	x"3010",	x"074e",	x"06b4",	
												x"0731",	x"0707",	x"0738",	x"06e3",	
												x"074c",	x"0725",	x"0762",	x"06f1",	
												x"0750",	x"0760",	x"0759",	x"072a",	
												x"0759",	x"072c",	x"079a",	x"0755",	
												x"079d",	x"0776",	x"076e",	x"0772",	
												x"079e",	x"0769",	x"0794",	x"075f",	
												x"0773",	x"0773",	x"076c",	x"0766",	
												x"0753",	x"0746",	x"0785",	x"0745",	
												x"0780",	x"0771",	x"07a7",	x"0771",	
												x"07af",	x"0776",	x"07ba",	x"0794",	
												x"07b8",	x"078a",	x"07b1",	x"07a8",	
												x"07a0",	x"0772",	x"07ce",	x"0778",	
												x"07b3",	x"0791",	x"0795",	x"077f",	
												x"079f",	x"0777",	x"07ec",	x"0761",	
												x"07ca",	x"078b",	x"07bf",	x"0797",	
												x"0759",	x"078b",	x"602f",	x"3010",	
												x"076e",	x"0717",	x"076f",	x"073c",	
												x"0758",	x"071e",	x"0738",	x"0701",	
												x"073b",	x"0715",	x"0769",	x"0740",	
												x"075c",	x"071f",	x"0769",	x"0737",	
												x"07c7",	x"0745",	x"07a2",	x"075d",	
												x"07ac",	x"0795",	x"07bc",	x"079c",	
												x"07a3",	x"0791",	x"07b3",	x"0799",	
												x"07c7",	x"0784",	x"0781",	x"078d",	
												x"07c9",	x"076f",	x"07d3",	x"07a7",	
												x"07dc",	x"0788",	x"07ef",	x"07b2",	
												x"080a",	x"07ac",	x"07de",	x"07bc",	
												x"07ff",	x"07ac",	x"07b7",	x"07ae",	
												x"07e6",	x"07a9",	x"07d2",	x"07c0",	
												x"07ce",	x"07a8",	x"07f0",	x"07a6",	
												x"080f",	x"07bd",	x"0807",	x"07cc",	
												x"0807",	x"07c1",	x"074f",	x"079c",	
												x"702f",	x"3010",	x"079a",	x"0728",	
												x"0777",	x"0747",	x"07ab",	x"0744",	
												x"0770",	x"074a",	x"07b5",	x"076e",	
												x"07e6",	x"0784",	x"07b1",	x"0773",	
												x"07ac",	x"078b",	x"0812",	x"0783",	
												x"0811",	x"07be",	x"081c",	x"07cd",	
												x"0834",	x"07da",	x"0816",	x"07e6",	
												x"0846",	x"07f8",	x"0804",	x"080a",	
												x"07d2",	x"07e3",	x"0826",	x"07c4",	
												x"0830",	x"0806",	x"0831",	x"07ef",	
												x"085d",	x"081e",	x"0834",	x"07fa",	
												x"0880",	x"081a",	x"086a",	x"082d",	
												x"082a",	x"0820",	x"0846",	x"0837",	
												x"084e",	x"082c",	x"085c",	x"0826",	
												x"0884",	x"0835",	x"0881",	x"0814",	
												x"0888",	x"083e",	x"0882",	x"083b",	
												x"069f",	x"081f",	x"0004",	x"000a",	
												x"7114",	x"0058",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"0011",	
												x"069a",	x"06eb",	x"0695",	x"0682",	
												x"0698",	x"067a",	x"068f",	x"067d",	
												x"06c0",	x"0673",	x"06eb",	x"06c5",	
												x"06cb",	x"06f8",	x"0684",	x"06c4",	
												x"06e0",	x"06ae",	x"06d6",	x"06e0",	
												x"06c0",	x"06c4",	x"06dc",	x"06dc",	
												x"06dc",	x"06d2",	x"06df",	x"06f0",	
												x"06de",	x"06dc",	x"068d",	x"06d6",	
												x"06cd",	x"069a",	x"06eb",	x"070a",	
												x"06b8",	x"06d5",	x"06c4",	x"06de",	
												x"06dc",	x"06a4",	x"06ef",	x"06e1",	
												x"06c3",	x"06ec",	x"06bb",	x"06c8",	
												x"06da",	x"06c5",	x"06e8",	x"06e7",	
												x"06f3",	x"06d8",	x"06f7",	x"06f6",	
												x"06d2",	x"06d7",	x"06da",	x"06c0",	
												x"06fd",	x"06c2",	x"06a6",	x"06f2",	
												x"1030",	x"0011",	x"0667",	x"06b4",	
												x"06a5",	x"0690",	x"0673",	x"06b7",	
												x"06a5",	x"0699",	x"06a3",	x"069f",	
												x"06c9",	x"06a6",	x"0696",	x"06c5",	
												x"06b0",	x"06c4",	x"06b4",	x"06a0",	
												x"06bf",	x"06bc",	x"06bc",	x"06e4",	
												x"06c0",	x"06ef",	x"06ba",	x"06d6",	
												x"06c2",	x"06cd",	x"06df",	x"06db",	
												x"067e",	x"06d0",	x"06b9",	x"069a",	
												x"06de",	x"06c1",	x"06ca",	x"06e2",	
												x"06c4",	x"06d0",	x"06c2",	x"06cf",	
												x"06d2",	x"06df",	x"06d0",	x"06e1",	
												x"06b6",	x"06d1",	x"06cb",	x"06c1",	
												x"06db",	x"06bd",	x"06fa",	x"06dd",	
												x"06fd",	x"0707",	x"06eb",	x"06ea",	
												x"06f9",	x"06da",	x"06ee",	x"0709",	
												x"0676",	x"06f9",	x"2030",	x"0011",	
												x"0673",	x"06ba",	x"069c",	x"0693",	
												x"066c",	x"067d",	x"068a",	x"0687",	
												x"068e",	x"06a3",	x"069f",	x"06b2",	
												x"0699",	x"06a5",	x"0686",	x"06c1",	
												x"06d2",	x"06ca",	x"06d1",	x"06df",	
												x"06d2",	x"06db",	x"06bc",	x"06d8",	
												x"06ba",	x"06b7",	x"06cd",	x"06bf",	
												x"06ab",	x"06be",	x"0687",	x"06ac",	
												x"06f0",	x"06a6",	x"06c8",	x"06c7",	
												x"06be",	x"06d0",	x"06ba",	x"06cd",	
												x"06e4",	x"06b3",	x"06d9",	x"06c2",	
												x"06d5",	x"06d4",	x"069d",	x"06cc",	
												x"06d9",	x"06ab",	x"06da",	x"06ce",	
												x"06cd",	x"06c8",	x"06d3",	x"06d5",	
												x"06eb",	x"06cf",	x"06e8",	x"06ee",	
												x"06e0",	x"06d4",	x"066d",	x"06be",	
												x"3030",	x"0011",	x"0676",	x"0675",	
												x"0690",	x"065f",	x"06ad",	x"0692",	
												x"068b",	x"0682",	x"06a6",	x"0688",	
												x"06ba",	x"06a5",	x"06b2",	x"069b",	
												x"068f",	x"0695",	x"06d7",	x"0699",	
												x"06b3",	x"06c5",	x"06b6",	x"06a0",	
												x"06b9",	x"06a8",	x"06c9",	x"06a1",	
												x"06b2",	x"06b1",	x"06c6",	x"0695",	
												x"0689",	x"06b6",	x"06c6",	x"06a4",	
												x"06cf",	x"06b6",	x"06cf",	x"06a0",	
												x"06f5",	x"06d7",	x"06f7",	x"06d1",	
												x"06d5",	x"06cb",	x"06cf",	x"06b3",	
												x"0696",	x"06cc",	x"06e4",	x"06aa",	
												x"070f",	x"06d5",	x"06f2",	x"06d7",	
												x"06de",	x"06dc",	x"0700",	x"06be",	
												x"06ec",	x"06ca",	x"0707",	x"06d1",	
												x"0699",	x"06e0",	x"0004",	x"000a",	
												x"0026",	x"e4a1",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"0012",	
												x"06af",	x"068f",	x"06a4",	x"06ad",	
												x"069a",	x"0692",	x"06d1",	x"069f",	
												x"06cf",	x"06b3",	x"06d0",	x"06ae",	
												x"06b9",	x"06ec",	x"06b8",	x"06a9",	
												x"06f0",	x"06c1",	x"06f9",	x"06e1",	
												x"06fd",	x"06ce",	x"0710",	x"06f2",	
												x"06e8",	x"06e0",	x"06e9",	x"06ec",	
												x"06ff",	x"06f0",	x"06d4",	x"06f0",	
												x"070c",	x"06e1",	x"071d",	x"0710",	
												x"070e",	x"0708",	x"0717",	x"0700",	
												x"071a",	x"06fa",	x"0715",	x"071c",	
												x"070a",	x"070f",	x"0709",	x"06f7",	
												x"0727",	x"0713",	x"0729",	x"071f",	
												x"0740",	x"0716",	x"0744",	x"0735",	
												x"0743",	x"0713",	x"0751",	x"071b",	
												x"0746",	x"0709",	x"06d0",	x"0719",	
												x"5030",	x"0012",	x"06dc",	x"06ee",	
												x"0700",	x"06bf",	x"06e0",	x"06f5",	
												x"06f7",	x"06e0",	x"0717",	x"06ea",	
												x"072b",	x"06e5",	x"073c",	x"0709",	
												x"0714",	x"0725",	x"0738",	x"06fa",	
												x"073c",	x"0719",	x"0749",	x"071a",	
												x"0744",	x"0736",	x"0739",	x"071a",	
												x"0734",	x"070f",	x"0725",	x"06f5",	
												x"0726",	x"0700",	x"0752",	x"06ff",	
												x"072c",	x"0729",	x"073a",	x"0703",	
												x"0743",	x"0717",	x"074f",	x"071b",	
												x"074f",	x"073b",	x"0760",	x"071c",	
												x"0751",	x"073d",	x"0764",	x"0705",	
												x"076f",	x"0740",	x"076d",	x"0742",	
												x"0781",	x"0730",	x"0780",	x"0730",	
												x"0775",	x"073c",	x"0769",	x"071e",	
												x"0704",	x"0731",	x"6030",	x"0012",	
												x"0725",	x"06f6",	x"0713",	x"06f7",	
												x"0739",	x"06c3",	x"0723",	x"06f3",	
												x"0736",	x"06f4",	x"0747",	x"0712",	
												x"074d",	x"0708",	x"0736",	x"072a",	
												x"076d",	x"071a",	x"0773",	x"0733",	
												x"0765",	x"0758",	x"0761",	x"074d",	
												x"0757",	x"0751",	x"0789",	x"0773",	
												x"075e",	x"0757",	x"075f",	x"073b",	
												x"075b",	x"073f",	x"077a",	x"076b",	
												x"077c",	x"0756",	x"077f",	x"0772",	
												x"076f",	x"0748",	x"0787",	x"074a",	
												x"0780",	x"0744",	x"077f",	x"0758",	
												x"078e",	x"0756",	x"07ac",	x"0775",	
												x"07a1",	x"077c",	x"07bf",	x"0784",	
												x"07bc",	x"0770",	x"07af",	x"0778",	
												x"07b3",	x"076f",	x"0760",	x"077c",	
												x"7030",	x"0012",	x"076e",	x"075d",	
												x"075b",	x"0727",	x"0771",	x"0713",	
												x"07ae",	x"073c",	x"0779",	x"0744",	
												x"0793",	x"0767",	x"079a",	x"0785",	
												x"0795",	x"076d",	x"07c0",	x"0768",	
												x"07c1",	x"07ab",	x"07c4",	x"07a6",	
												x"07ca",	x"0795",	x"07bc",	x"07a8",	
												x"07ce",	x"079b",	x"07c9",	x"07af",	
												x"07c6",	x"07ac",	x"07f9",	x"07b9",	
												x"07ee",	x"07c1",	x"0812",	x"07c2",	
												x"07fc",	x"07d9",	x"07e0",	x"07db",	
												x"07f9",	x"07cb",	x"07e3",	x"07cc",	
												x"07e9",	x"07ef",	x"07ff",	x"07d4",	
												x"081b",	x"07ed",	x"0810",	x"07e7",	
												x"0852",	x"0801",	x"0836",	x"0811",	
												x"0835",	x"0819",	x"0822",	x"081d",	
												x"064f",	x"07fe",	x"0004",	x"000a",	
												x"4d6e",	x"220f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"1013",	
												x"0646",	x"0647",	x"0654",	x"065c",	
												x"065c",	x"065f",	x"067b",	x"066b",	
												x"0683",	x"06a1",	x"0683",	x"066d",	
												x"0675",	x"065e",	x"0667",	x"0667",	
												x"067f",	x"0677",	x"0674",	x"06c1",	
												x"06a2",	x"0678",	x"0691",	x"0696",	
												x"069c",	x"0696",	x"069d",	x"06ba",	
												x"0695",	x"06a3",	x"0652",	x"06ad",	
												x"066f",	x"066e",	x"0689",	x"065e",	
												x"0678",	x"0676",	x"067e",	x"0685",	
												x"0695",	x"0695",	x"06ba",	x"067e",	
												x"068e",	x"06b2",	x"0642",	x"06a6",	
												x"067d",	x"0655",	x"06a7",	x"0695",	
												x"06a3",	x"069b",	x"068e",	x"06b8",	
												x"068f",	x"069b",	x"0698",	x"06a0",	
												x"0694",	x"067a",	x"061e",	x"067e",	
												x"1030",	x"1013",	x"062d",	x"0633",	
												x"0641",	x"0632",	x"064c",	x"063f",	
												x"0671",	x"066b",	x"066d",	x"0672",	
												x"0693",	x"066f",	x"0665",	x"068a",	
												x"065a",	x"068c",	x"0663",	x"066e",	
												x"0679",	x"0683",	x"0686",	x"067a",	
												x"0691",	x"06aa",	x"0681",	x"0680",	
												x"068b",	x"0698",	x"067f",	x"068a",	
												x"0667",	x"0692",	x"0658",	x"0665",	
												x"0663",	x"066d",	x"068a",	x"0672",	
												x"0674",	x"069a",	x"0698",	x"067c",	
												x"06aa",	x"06b2",	x"068e",	x"06bb",	
												x"0683",	x"068f",	x"0677",	x"067d",	
												x"0695",	x"0682",	x"06c3",	x"06aa",	
												x"0698",	x"06b2",	x"06ac",	x"06a2",	
												x"068d",	x"0692",	x"0698",	x"0693",	
												x"064e",	x"06a3",	x"2030",	x"1013",	
												x"063b",	x"066a",	x"064e",	x"0650",	
												x"065b",	x"0652",	x"063a",	x"0658",	
												x"065b",	x"065b",	x"067a",	x"066b",	
												x"0647",	x"0663",	x"063e",	x"0664",	
												x"0673",	x"0681",	x"0669",	x"0687",	
												x"0649",	x"066e",	x"067d",	x"0666",	
												x"0680",	x"067c",	x"067e",	x"0673",	
												x"0672",	x"067f",	x"0646",	x"0678",	
												x"0685",	x"0644",	x"0674",	x"066a",	
												x"0660",	x"064e",	x"0672",	x"0675",	
												x"0699",	x"067c",	x"069e",	x"0696",	
												x"067a",	x"068d",	x"064d",	x"0668",	
												x"068a",	x"0667",	x"0698",	x"0689",	
												x"068f",	x"066d",	x"0693",	x"0691",	
												x"068a",	x"067a",	x"0678",	x"0677",	
												x"0685",	x"0663",	x"063e",	x"066e",	
												x"3030",	x"1013",	x"0634",	x"063c",	
												x"063f",	x"0617",	x"065b",	x"0629",	
												x"0656",	x"0643",	x"0661",	x"064f",	
												x"0656",	x"0657",	x"0675",	x"0655",	
												x"064a",	x"066d",	x"0658",	x"0638",	
												x"0652",	x"0662",	x"066c",	x"0657",	
												x"067c",	x"0665",	x"066d",	x"0656",	
												x"0676",	x"0670",	x"0666",	x"0665",	
												x"0663",	x"064e",	x"0663",	x"065e",	
												x"066e",	x"066e",	x"0676",	x"0677",	
												x"0677",	x"067e",	x"067e",	x"0674",	
												x"0677",	x"066c",	x"068c",	x"0670",	
												x"0686",	x"066c",	x"069e",	x"0664",	
												x"0693",	x"0674",	x"0699",	x"0678",	
												x"069e",	x"068f",	x"0696",	x"067f",	
												x"0695",	x"0689",	x"0689",	x"0666",	
												x"064c",	x"066d",	x"0004",	x"000a",	
												x"da78",	x"ff74",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"1014",	
												x"064f",	x"062b",	x"066c",	x"061e",	
												x"0683",	x"0640",	x"0689",	x"065d",	
												x"0681",	x"0662",	x"0686",	x"0683",	
												x"0692",	x"067d",	x"067b",	x"0684",	
												x"06a1",	x"0673",	x"0694",	x"0688",	
												x"068e",	x"067d",	x"0699",	x"0692",	
												x"06a9",	x"0692",	x"06a2",	x"06a1",	
												x"0698",	x"06a7",	x"067a",	x"06a0",	
												x"06ae",	x"0689",	x"06af",	x"06b4",	
												x"069b",	x"06a0",	x"06ad",	x"06ba",	
												x"06a2",	x"06bf",	x"06c8",	x"06ac",	
												x"06ca",	x"06b5",	x"06af",	x"06bc",	
												x"06c2",	x"06ab",	x"06cc",	x"06a8",	
												x"06c6",	x"06ca",	x"06d6",	x"06d8",	
												x"06e0",	x"06be",	x"06cc",	x"06c5",	
												x"06df",	x"069b",	x"0698",	x"06bb",	
												x"5030",	x"1014",	x"0680",	x"0696",	
												x"06a3",	x"0669",	x"06a2",	x"0673",	
												x"06b2",	x"06ad",	x"06cf",	x"06a6",	
												x"06d7",	x"06b1",	x"06cd",	x"06cb",	
												x"06bc",	x"06de",	x"06ce",	x"06c3",	
												x"06cf",	x"06c1",	x"06db",	x"06c5",	
												x"06de",	x"06d6",	x"06c9",	x"06bc",	
												x"06c9",	x"06b0",	x"06ce",	x"06b3",	
												x"06b7",	x"06be",	x"06ce",	x"06b3",	
												x"06de",	x"06c4",	x"06e8",	x"06cb",	
												x"06fe",	x"06d1",	x"06f0",	x"06db",	
												x"06f8",	x"06db",	x"06fd",	x"06e5",	
												x"06f0",	x"06df",	x"06f6",	x"06cb",	
												x"0712",	x"06c4",	x"070b",	x"06cb",	
												x"06f8",	x"06e8",	x"06ec",	x"06ce",	
												x"0708",	x"06df",	x"06fb",	x"06e4",	
												x"06a8",	x"06e6",	x"6030",	x"1014",	
												x"06bd",	x"067e",	x"06cf",	x"0682",	
												x"06b4",	x"0681",	x"06d0",	x"06ad",	
												x"06db",	x"06df",	x"06f8",	x"06cb",	
												x"06f5",	x"06c7",	x"06bc",	x"06dc",	
												x"06fc",	x"06c1",	x"070a",	x"06e4",	
												x"0715",	x"06c3",	x"070c",	x"06fc",	
												x"0704",	x"06f2",	x"06ff",	x"06f1",	
												x"0721",	x"06db",	x"06d3",	x"06da",	
												x"0711",	x"06c9",	x"06f9",	x"0702",	
												x"070b",	x"06e6",	x"072f",	x"070b",	
												x"0728",	x"0723",	x"072a",	x"071a",	
												x"071d",	x"070a",	x"0706",	x"0701",	
												x"073a",	x"06f7",	x"0731",	x"0726",	
												x"072d",	x"0710",	x"072d",	x"0704",	
												x"0740",	x"0716",	x"0746",	x"0725",	
												x"072a",	x"071d",	x"070b",	x"0707",	
												x"7030",	x"1014",	x"0712",	x"06d9",	
												x"0706",	x"06e3",	x"072a",	x"06f5",	
												x"0729",	x"071d",	x"0711",	x"06ff",	
												x"0722",	x"0713",	x"071b",	x"06fa",	
												x"0736",	x"071a",	x"0762",	x"072a",	
												x"0745",	x"074b",	x"0757",	x"072b",	
												x"0770",	x"075b",	x"0775",	x"0744",	
												x"077c",	x"075a",	x"0761",	x"0757",	
												x"0762",	x"0752",	x"076e",	x"0738",	
												x"0772",	x"0758",	x"0772",	x"0768",	
												x"07b5",	x"0762",	x"07b9",	x"077f",	
												x"0799",	x"0789",	x"0776",	x"0759",	
												x"075a",	x"0759",	x"07a1",	x"075a",	
												x"0792",	x"079b",	x"078b",	x"07a8",	
												x"07c1",	x"0790",	x"07bc",	x"0790",	
												x"07b7",	x"07b7",	x"07a8",	x"079a",	
												x"0709",	x"0782",	x"0004",	x"000a",	
												x"1ce9",	x"3617",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"2015",	
												x"0701",	x"0749",	x"0702",	x"0703",	
												x"070f",	x"070c",	x"0720",	x"0719",	
												x"074d",	x"072c",	x"074e",	x"073f",	
												x"074f",	x"0743",	x"072d",	x"076a",	
												x"0729",	x"073c",	x"0724",	x"0762",	
												x"0751",	x"074e",	x"0758",	x"075a",	
												x"0769",	x"0774",	x"0773",	x"0792",	
												x"074e",	x"0782",	x"06f3",	x"0757",	
												x"0734",	x"0741",	x"0755",	x"074b",	
												x"0734",	x"0753",	x"0752",	x"0749",	
												x"0741",	x"0753",	x"0747",	x"0755",	
												x"0746",	x"0753",	x"071c",	x"075b",	
												x"0732",	x"071f",	x"074c",	x"0734",	
												x"074f",	x"0742",	x"076a",	x"0751",	
												x"073c",	x"071f",	x"077d",	x"0745",	
												x"076f",	x"0744",	x"06e1",	x"0753",	
												x"1030",	x"2015",	x"06f6",	x"06ed",	
												x"0705",	x"0706",	x"06fd",	x"0701",	
												x"0740",	x"06f2",	x"072c",	x"0731",	
												x"0731",	x"073d",	x"072c",	x"073d",	
												x"070c",	x"074b",	x"0733",	x"0716",	
												x"0734",	x"0741",	x"0770",	x"0731",	
												x"0790",	x"0785",	x"075d",	x"0752",	
												x"075d",	x"0770",	x"0747",	x"0744",	
												x"0706",	x"0746",	x"0725",	x"071d",	
												x"0749",	x"074f",	x"0757",	x"075a",	
												x"073e",	x"075c",	x"072e",	x"0737",	
												x"077c",	x"0740",	x"0769",	x"0764",	
												x"0720",	x"0757",	x"075a",	x"0736",	
												x"076a",	x"075f",	x"0763",	x"0766",	
												x"0752",	x"0765",	x"0745",	x"074c",	
												x"0789",	x"074c",	x"0763",	x"0771",	
												x"06eb",	x"0762",	x"2030",	x"2015",	
												x"070b",	x"06ec",	x"06fc",	x"0712",	
												x"0708",	x"070d",	x"0713",	x"0742",	
												x"071f",	x"072d",	x"0720",	x"0743",	
												x"0711",	x"0732",	x"06f5",	x"072c",	
												x"0705",	x"070f",	x"0709",	x"0740",	
												x"0724",	x"0736",	x"0756",	x"0730",	
												x"074a",	x"0758",	x"0734",	x"074f",	
												x"0759",	x"0752",	x"06c4",	x"0734",	
												x"0727",	x"071c",	x"071b",	x"0728",	
												x"0727",	x"070e",	x"0727",	x"0736",	
												x"072c",	x"0731",	x"0767",	x"0743",	
												x"073c",	x"074c",	x"071f",	x"073f",	
												x"0747",	x"0731",	x"0752",	x"073d",	
												x"073e",	x"0726",	x"074b",	x"0762",	
												x"074b",	x"0740",	x"0747",	x"0732",	
												x"0737",	x"0731",	x"06d2",	x"0752",	
												x"3030",	x"2015",	x"06e7",	x"06cf",	
												x"06f1",	x"06ce",	x"06f1",	x"0700",	
												x"06f6",	x"0705",	x"0712",	x"06fe",	
												x"072e",	x"0708",	x"0708",	x"0718",	
												x"06ec",	x"0719",	x"0709",	x"0704",	
												x"072d",	x"0722",	x"0749",	x"073c",	
												x"0738",	x"0736",	x"073f",	x"0727",	
												x"073a",	x"0751",	x"072e",	x"0715",	
												x"06f2",	x"0733",	x"072c",	x"0707",	
												x"0730",	x"072a",	x"0739",	x"073b",	
												x"074d",	x"0738",	x"074e",	x"0740",	
												x"0750",	x"073d",	x"074d",	x"073a",	
												x"0703",	x"0741",	x"0734",	x"0713",	
												x"0756",	x"072c",	x"0768",	x"0732",	
												x"0762",	x"0732",	x"075c",	x"0738",	
												x"077b",	x"074f",	x"0774",	x"0738",	
												x"070a",	x"0742",	x"0004",	x"000a",	
												x"39b8",	x"a084",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"2016",	
												x"0711",	x"070a",	x"0714",	x"0724",	
												x"0742",	x"071e",	x"074a",	x"071e",	
												x"074a",	x"0730",	x"0749",	x"0761",	
												x"0741",	x"0733",	x"0728",	x"0744",	
												x"0736",	x"074c",	x"0761",	x"0750",	
												x"075d",	x"076e",	x"0774",	x"0760",	
												x"0783",	x"0758",	x"077e",	x"077e",	
												x"0761",	x"074d",	x"0737",	x"074b",	
												x"076b",	x"0756",	x"0769",	x"075d",	
												x"0778",	x"076e",	x"0794",	x"077f",	
												x"077e",	x"077a",	x"078d",	x"077e",	
												x"0780",	x"079b",	x"078d",	x"077f",	
												x"0792",	x"077c",	x"0787",	x"0791",	
												x"079e",	x"077e",	x"07ba",	x"0799",	
												x"07a5",	x"079a",	x"079e",	x"0799",	
												x"07c4",	x"0792",	x"0730",	x"07a9",	
												x"5030",	x"2016",	x"074f",	x"0748",	
												x"0775",	x"0723",	x"076d",	x"074e",	
												x"0775",	x"0764",	x"079a",	x"0773",	
												x"0775",	x"0773",	x"0773",	x"077e",	
												x"07a0",	x"075b",	x"07a8",	x"07a5",	
												x"07ad",	x"07a4",	x"079d",	x"0791",	
												x"07d0",	x"0799",	x"07af",	x"07b5",	
												x"07ad",	x"07a8",	x"07bc",	x"07aa",	
												x"0792",	x"0784",	x"07ae",	x"0765",	
												x"07bb",	x"07aa",	x"07d9",	x"079d",	
												x"07c7",	x"07b0",	x"07bb",	x"07a7",	
												x"07df",	x"07aa",	x"07d3",	x"07ac",	
												x"07b5",	x"07a5",	x"07bb",	x"0794",	
												x"07da",	x"07a4",	x"07e0",	x"07a2",	
												x"07fb",	x"07a1",	x"07f7",	x"07ac",	
												x"07ec",	x"07b5",	x"07de",	x"07af",	
												x"0778",	x"07af",	x"6030",	x"2016",	
												x"0777",	x"0751",	x"076d",	x"075d",	
												x"0771",	x"0759",	x"079c",	x"0757",	
												x"079e",	x"0779",	x"07ae",	x"077c",	
												x"07a9",	x"0788",	x"07c1",	x"0793",	
												x"07e2",	x"0783",	x"07e7",	x"078d",	
												x"07e5",	x"07c3",	x"07ff",	x"07c1",	
												x"07ed",	x"07b7",	x"07f8",	x"07ce",	
												x"07cd",	x"07aa",	x"07db",	x"07c6",	
												x"07e2",	x"07bf",	x"07d8",	x"07df",	
												x"0804",	x"07c0",	x"07fe",	x"07e3",	
												x"07f8",	x"07be",	x"0802",	x"0803",	
												x"080c",	x"07c3",	x"0800",	x"07f9",	
												x"0804",	x"07ef",	x"081a",	x"07df",	
												x"0827",	x"07de",	x"081d",	x"0804",	
												x"0815",	x"07f8",	x"081f",	x"07d7",	
												x"0835",	x"07e8",	x"07e0",	x"07f1",	
												x"7030",	x"2016",	x"07bb",	x"07a4",	
												x"07fb",	x"07a8",	x"07e4",	x"077e",	
												x"0819",	x"07c7",	x"0809",	x"07e8",	
												x"081c",	x"0815",	x"0810",	x"0817",	
												x"07e7",	x"07ed",	x"0838",	x"07e7",	
												x"083f",	x"0822",	x"0849",	x"0833",	
												x"0896",	x"084a",	x"0863",	x"0825",	
												x"0855",	x"082a",	x"0855",	x"0833",	
												x"0840",	x"081c",	x"0843",	x"0837",	
												x"088d",	x"083f",	x"0880",	x"0838",	
												x"0880",	x"086d",	x"0874",	x"0857",	
												x"087f",	x"084e",	x"088a",	x"0858",	
												x"0867",	x"0856",	x"0885",	x"084d",	
												x"088e",	x"087c",	x"08a0",	x"088c",	
												x"0893",	x"0890",	x"08af",	x"087c",	
												x"08bd",	x"0898",	x"0894",	x"088f",	
												x"0710",	x"0896",	x"0004",	x"000a",	
												x"88bc",	x"e037",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"3017",	
												x"06d2",	x"06f3",	x"06d2",	x"06dd",	
												x"06d4",	x"06d0",	x"06c9",	x"06ec",	
												x"06ee",	x"0709",	x"0713",	x"06f7",	
												x"0717",	x"0733",	x"06f2",	x"071f",	
												x"0723",	x"06fa",	x"071c",	x"0729",	
												x"0717",	x"071f",	x"0743",	x"0755",	
												x"073a",	x"070d",	x"073e",	x"0726",	
												x"06f7",	x"0749",	x"06d4",	x"06fe",	
												x"070f",	x"06fc",	x"0717",	x"0717",	
												x"06f5",	x"0713",	x"072f",	x"0702",	
												x"0717",	x"06fe",	x"0766",	x"073b",	
												x"0737",	x"0755",	x"06f3",	x"071e",	
												x"0710",	x"06e7",	x"0716",	x"0717",	
												x"0722",	x"0715",	x"0727",	x"073b",	
												x"072c",	x"0710",	x"0765",	x"0727",	
												x"0750",	x"073f",	x"06cf",	x"071c",	
												x"1030",	x"3017",	x"06d9",	x"06ea",	
												x"06fa",	x"06eb",	x"06dc",	x"06f0",	
												x"06e1",	x"06d7",	x"06ec",	x"06df",	
												x"0719",	x"0719",	x"06e4",	x"0716",	
												x"06d8",	x"06f2",	x"070d",	x"06f2",	
												x"0729",	x"0733",	x"0712",	x"073c",	
												x"0718",	x"0743",	x"071e",	x"070a",	
												x"070b",	x"0718",	x"070f",	x"0719",	
												x"06dc",	x"0736",	x"0702",	x"06d1",	
												x"06e8",	x"0722",	x"0705",	x"06ee",	
												x"0718",	x"0742",	x"0707",	x"0724",	
												x"0729",	x"073d",	x"0730",	x"072e",	
												x"06fe",	x"071c",	x"06f6",	x"06f1",	
												x"06fb",	x"06fa",	x"0721",	x"0719",	
												x"072a",	x"0719",	x"0740",	x"0715",	
												x"0739",	x"073c",	x"0734",	x"072e",	
												x"06ed",	x"072c",	x"2030",	x"3017",	
												x"06e6",	x"06ee",	x"06eb",	x"06f4",	
												x"06c8",	x"06e6",	x"06d0",	x"06da",	
												x"06d6",	x"0701",	x"06fc",	x"06f9",	
												x"06ee",	x"0704",	x"06ef",	x"071a",	
												x"070b",	x"0712",	x"06f8",	x"0727",	
												x"0712",	x"0737",	x"070b",	x"0705",	
												x"0706",	x"070a",	x"0723",	x"0718",	
												x"06f7",	x"06f8",	x"06e7",	x"0704",	
												x"06ec",	x"06f7",	x"06ed",	x"06f3",	
												x"06ec",	x"06d3",	x"06f6",	x"06f2",	
												x"072d",	x"0706",	x"072e",	x"0734",	
												x"071f",	x"0727",	x"06f2",	x"070a",	
												x"06f5",	x"06f8",	x"06f9",	x"06f3",	
												x"0708",	x"06fe",	x"071c",	x"0705",	
												x"072f",	x"070e",	x"0717",	x"071d",	
												x"0730",	x"06f7",	x"06d5",	x"0712",	
												x"3030",	x"3017",	x"06dc",	x"06d2",	
												x"06e1",	x"06e5",	x"06b1",	x"06d2",	
												x"06db",	x"06c9",	x"06e7",	x"06b6",	
												x"06e6",	x"06dc",	x"06ec",	x"06e5",	
												x"06de",	x"06d3",	x"06e4",	x"06e3",	
												x"06ff",	x"0712",	x"0722",	x"06fd",	
												x"06ee",	x"071c",	x"0701",	x"06e2",	
												x"06f7",	x"06f6",	x"06f1",	x"06f8",	
												x"06d0",	x"06e5",	x"06f7",	x"06cd",	
												x"0706",	x"06f8",	x"0711",	x"06ef",	
												x"06f4",	x"0711",	x"0716",	x"06e2",	
												x"0728",	x"0718",	x"0715",	x"0708",	
												x"06fe",	x"06ee",	x"071d",	x"06fa",	
												x"070f",	x"0727",	x"0717",	x"06fe",	
												x"0737",	x"0707",	x"0731",	x"0710",	
												x"0746",	x"071c",	x"0715",	x"06fa",	
												x"06e5",	x"0708",	x"0004",	x"000a",	
												x"2260",	x"c826",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"3018",	
												x"06f1",	x"06ce",	x"06f9",	x"06d2",	
												x"0709",	x"06fd",	x"06ec",	x"06fb",	
												x"0704",	x"06e8",	x"070a",	x"0708",	
												x"070a",	x"071b",	x"070f",	x"0704",	
												x"070e",	x"0717",	x"071a",	x"072b",	
												x"072a",	x"0711",	x"072e",	x"070f",	
												x"072f",	x"0718",	x"073e",	x"072a",	
												x"0729",	x"073c",	x"0715",	x"072b",	
												x"0729",	x"0729",	x"072d",	x"0721",	
												x"072b",	x"0728",	x"073e",	x"0735",	
												x"0751",	x"0736",	x"0757",	x"0737",	
												x"075f",	x"073d",	x"0710",	x"0758",	
												x"0743",	x"072f",	x"0752",	x"0740",	
												x"075c",	x"074e",	x"0788",	x"0769",	
												x"0781",	x"0767",	x"0775",	x"0771",	
												x"0769",	x"074a",	x"074b",	x"0742",	
												x"5030",	x"3018",	x"070f",	x"0735",	
												x"0730",	x"06f9",	x"072a",	x"06ef",	
												x"0741",	x"0726",	x"0757",	x"0722",	
												x"0755",	x"074f",	x"0755",	x"073b",	
												x"0761",	x"073b",	x"075e",	x"0756",	
												x"075c",	x"0764",	x"075a",	x"0766",	
												x"0755",	x"0765",	x"0783",	x"0755",	
												x"0766",	x"076a",	x"0764",	x"076a",	
												x"0760",	x"075d",	x"0756",	x"072a",	
												x"075c",	x"0748",	x"0773",	x"075f",	
												x"078b",	x"0770",	x"07bb",	x"0774",	
												x"07a7",	x"078f",	x"078e",	x"078e",	
												x"0779",	x"0778",	x"0793",	x"0757",	
												x"0783",	x"0747",	x"07ae",	x"0778",	
												x"07ac",	x"0782",	x"07be",	x"077b",	
												x"07bf",	x"0783",	x"079e",	x"078f",	
												x"0755",	x"0776",	x"6030",	x"3018",	
												x"0767",	x"0723",	x"074f",	x"0751",	
												x"0742",	x"0730",	x"0770",	x"0731",	
												x"076e",	x"0774",	x"075c",	x"075d",	
												x"0761",	x"0749",	x"0773",	x"075b",	
												x"078e",	x"076a",	x"0798",	x"0779",	
												x"079c",	x"078f",	x"07a9",	x"0797",	
												x"079b",	x"078f",	x"0799",	x"079c",	
												x"07a0",	x"0774",	x"076f",	x"0774",	
												x"078f",	x"0779",	x"07ad",	x"0793",	
												x"07ac",	x"0791",	x"07c7",	x"078b",	
												x"07c0",	x"079c",	x"07d2",	x"07b3",	
												x"07c4",	x"07b1",	x"07c4",	x"07b0",	
												x"07d1",	x"07a7",	x"07aa",	x"07a5",	
												x"07cf",	x"079c",	x"07ff",	x"07b4",	
												x"07da",	x"07c2",	x"07e5",	x"07c9",	
												x"07e0",	x"07a4",	x"0760",	x"07bc",	
												x"7030",	x"3018",	x"07a3",	x"075c",	
												x"07a7",	x"0783",	x"07a4",	x"077f",	
												x"07b2",	x"077f",	x"07c4",	x"079c",	
												x"07e4",	x"07bc",	x"07a4",	x"07ba",	
												x"07b3",	x"07c1",	x"0814",	x"07da",	
												x"07f5",	x"07f8",	x"07f3",	x"07f6",	
												x"080d",	x"07f3",	x"082d",	x"0805",	
												x"0838",	x"081e",	x"080d",	x"0807",	
												x"07cf",	x"07fc",	x"080e",	x"07cf",	
												x"081e",	x"07fb",	x"081c",	x"080c",	
												x"0850",	x"081f",	x"0838",	x"081f",	
												x"085f",	x"085a",	x"0836",	x"0854",	
												x"0826",	x"0845",	x"0832",	x"0847",	
												x"0863",	x"0846",	x"0866",	x"083f",	
												x"0874",	x"0850",	x"0892",	x"0848",	
												x"0885",	x"085a",	x"0863",	x"0864",	
												x"06b6",	x"0867",	x"0004",	x"000a",	
												x"68b9",	x"0535",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"0019",	
												x"06c1",	x"06dc",	x"06c2",	x"06c2",	
												x"06d8",	x"06c8",	x"06ce",	x"06cf",	
												x"06b9",	x"06ae",	x"0692",	x"069b",	
												x"069f",	x"0684",	x"0670",	x"06a5",	
												x"06b4",	x"067e",	x"06ad",	x"06b6",	
												x"06b9",	x"06ab",	x"06c5",	x"06be",	
												x"06bf",	x"06c1",	x"06cc",	x"06e3",	
												x"06d1",	x"06d4",	x"06a2",	x"06ba",	
												x"06e0",	x"06bb",	x"06c3",	x"06c7",	
												x"06d3",	x"06c4",	x"06d0",	x"06e5",	
												x"06f2",	x"06a5",	x"0706",	x"06e5",	
												x"0708",	x"0715",	x"0693",	x"06ec",	
												x"06c3",	x"0692",	x"06c6",	x"06ca",	
												x"06d1",	x"06c9",	x"06de",	x"06dd",	
												x"06e2",	x"06aa",	x"0717",	x"06e7",	
												x"070b",	x"06ee",	x"06b3",	x"06df",	
												x"1031",	x"0019",	x"06a9",	x"06bc",	
												x"06ab",	x"06c8",	x"06a3",	x"0697",	
												x"06c0",	x"069f",	x"0682",	x"06ac",	
												x"0686",	x"0689",	x"069e",	x"0680",	
												x"066b",	x"067c",	x"068e",	x"067f",	
												x"0688",	x"0690",	x"06b1",	x"069b",	
												x"06d2",	x"06ae",	x"06f0",	x"06d4",	
												x"06d2",	x"06ef",	x"06e9",	x"06d6",	
												x"069c",	x"06cf",	x"06c4",	x"069f",	
												x"06b3",	x"06db",	x"06b3",	x"06c4",	
												x"06bf",	x"06d0",	x"06c4",	x"06d4",	
												x"06b9",	x"06c7",	x"06da",	x"06e0",	
												x"0694",	x"06d0",	x"06d9",	x"06b2",	
												x"06d1",	x"06c9",	x"06b9",	x"06c7",	
												x"06c2",	x"06ca",	x"06f2",	x"06ee",	
												x"06fc",	x"06ea",	x"06ff",	x"0703",	
												x"06b3",	x"06ee",	x"2031",	x"0019",	
												x"06ab",	x"06b5",	x"06af",	x"06aa",	
												x"06a0",	x"0688",	x"069a",	x"068e",	
												x"067f",	x"068c",	x"0696",	x"0695",	
												x"0679",	x"0698",	x"0632",	x"0687",	
												x"0699",	x"0667",	x"0697",	x"0694",	
												x"068f",	x"06ab",	x"06ad",	x"06b0",	
												x"06e0",	x"06b7",	x"06ec",	x"06ee",	
												x"06c0",	x"06b0",	x"068e",	x"06b8",	
												x"06c3",	x"06b0",	x"06b3",	x"06c9",	
												x"06b3",	x"06bc",	x"06d6",	x"06bd",	
												x"06cd",	x"06cf",	x"06d6",	x"06c8",	
												x"06ea",	x"06c9",	x"069e",	x"06cc",	
												x"06ca",	x"06c3",	x"06c8",	x"06a0",	
												x"06bf",	x"069e",	x"06c4",	x"06d1",	
												x"06ec",	x"06c9",	x"0700",	x"06d8",	
												x"0712",	x"06db",	x"0689",	x"06e0",	
												x"3031",	x"0019",	x"0688",	x"0677",	
												x"069b",	x"0673",	x"06b1",	x"068f",	
												x"06a9",	x"068f",	x"06bb",	x"067e",	
												x"06b2",	x"06a7",	x"0668",	x"068b",	
												x"065f",	x"0672",	x"068f",	x"065d",	
												x"06a2",	x"0680",	x"06ba",	x"06a1",	
												x"06f4",	x"06c2",	x"06f6",	x"06cc",	
												x"06d5",	x"06bd",	x"06d9",	x"06d3",	
												x"069c",	x"06d8",	x"06ad",	x"06c5",	
												x"06dd",	x"06ad",	x"06c1",	x"06d5",	
												x"06f4",	x"06c3",	x"06ea",	x"06b6",	
												x"06e9",	x"06c6",	x"06ef",	x"06d0",	
												x"06ab",	x"06cc",	x"06ee",	x"06a9",	
												x"06e8",	x"069a",	x"06ec",	x"06ab",	
												x"0705",	x"06db",	x"0741",	x"06dd",	
												x"071a",	x"06e5",	x"0729",	x"06dd",	
												x"06b5",	x"06f4",	x"0004",	x"000a",	
												x"0025",	x"e138",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"001a",	
												x"06cd",	x"06ac",	x"06da",	x"06a4",	
												x"06ce",	x"06b2",	x"06d9",	x"06b0",	
												x"06db",	x"06ba",	x"06b4",	x"0695",	
												x"06a2",	x"0697",	x"0691",	x"0694",	
												x"06dd",	x"0695",	x"06f4",	x"06cb",	
												x"0702",	x"06b5",	x"073e",	x"06d6",	
												x"0716",	x"06d9",	x"0714",	x"06ea",	
												x"0715",	x"0704",	x"06fa",	x"06f2",	
												x"0723",	x"06d3",	x"0723",	x"0727",	
												x"0735",	x"0717",	x"072d",	x"070e",	
												x"073b",	x"0705",	x"0742",	x"071b",	
												x"0739",	x"0727",	x"0720",	x"0704",	
												x"0736",	x"06fc",	x"072d",	x"0710",	
												x"0722",	x"070b",	x"0750",	x"071c",	
												x"078b",	x"072e",	x"0763",	x"0754",	
												x"0756",	x"0726",	x"0707",	x"0725",	
												x"5031",	x"001a",	x"0713",	x"0704",	
												x"0701",	x"06d5",	x"070b",	x"06bd",	
												x"0717",	x"06d4",	x"0713",	x"06c4",	
												x"072f",	x"06ed",	x"06f0",	x"06d4",	
												x"070c",	x"06c2",	x"0738",	x"06bc",	
												x"0745",	x"06fa",	x"075d",	x"070f",	
												x"0757",	x"0701",	x"0750",	x"0712",	
												x"0771",	x"0746",	x"0746",	x"0702",	
												x"0722",	x"0723",	x"0734",	x"070b",	
												x"0733",	x"0711",	x"0741",	x"0700",	
												x"076f",	x"0716",	x"0775",	x"0734",	
												x"0763",	x"0731",	x"0779",	x"0721",	
												x"076c",	x"0737",	x"077d",	x"071c",	
												x"0775",	x"073b",	x"0795",	x"0712",	
												x"07a1",	x"072d",	x"07e1",	x"072c",	
												x"0795",	x"075c",	x"077d",	x"0746",	
												x"06f6",	x"0738",	x"6031",	x"001a",	
												x"0712",	x"06e0",	x"0719",	x"06de",	
												x"0730",	x"06f7",	x"0722",	x"06fb",	
												x"0730",	x"06e2",	x"072b",	x"06f3",	
												x"0717",	x"06ca",	x"06d6",	x"06d1",	
												x"0765",	x"06bc",	x"0770",	x"0707",	
												x"0774",	x"0718",	x"0772",	x"073a",	
												x"0764",	x"074d",	x"0780",	x"0768",	
												x"078f",	x"0741",	x"075d",	x"073d",	
												x"077d",	x"0739",	x"0778",	x"0741",	
												x"07a3",	x"076a",	x"07a4",	x"0759",	
												x"079a",	x"0763",	x"0797",	x"0759",	
												x"07a3",	x"0753",	x"0777",	x"0763",	
												x"07a6",	x"0751",	x"07b2",	x"076c",	
												x"07ba",	x"0762",	x"07f4",	x"0780",	
												x"07d0",	x"0783",	x"07d4",	x"0792",	
												x"07d1",	x"0795",	x"0747",	x"0779",	
												x"7031",	x"001a",	x"074f",	x"072a",	
												x"0758",	x"0724",	x"0781",	x"071e",	
												x"078f",	x"075a",	x"077b",	x"074c",	
												x"077a",	x"073e",	x"078a",	x"0731",	
												x"072f",	x"0727",	x"07af",	x"0705",	
												x"07b9",	x"077d",	x"07ff",	x"076d",	
												x"0806",	x"0792",	x"07f4",	x"07ab",	
												x"07d6",	x"07c1",	x"0801",	x"07b6",	
												x"07c2",	x"07a8",	x"0800",	x"07ac",	
												x"080d",	x"07b6",	x"0810",	x"07ba",	
												x"0821",	x"07c4",	x"0819",	x"07d3",	
												x"0813",	x"07f9",	x"080b",	x"07bb",	
												x"07ce",	x"07cc",	x"07fd",	x"07bc",	
												x"0822",	x"07f0",	x"0833",	x"07e5",	
												x"0843",	x"0811",	x"0854",	x"0833",	
												x"0851",	x"0822",	x"0817",	x"0829",	
												x"066b",	x"07f8",	x"0004",	x"000a",	
												x"5442",	x"1e28",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"101b",	
												x"067a",	x"0667",	x"0682",	x"067e",	
												x"0659",	x"0666",	x"0654",	x"0661",	
												x"0638",	x"064f",	x"065e",	x"064d",	
												x"064d",	x"0643",	x"05ff",	x"0632",	
												x"0632",	x"0625",	x"0679",	x"0664",	
												x"0681",	x"0681",	x"06a2",	x"068c",	
												x"068f",	x"06b3",	x"0683",	x"06a4",	
												x"0677",	x"0696",	x"066c",	x"069d",	
												x"066b",	x"0680",	x"0659",	x"066e",	
												x"0664",	x"0677",	x"06ba",	x"066c",	
												x"068d",	x"0674",	x"0696",	x"068f",	
												x"069d",	x"06a2",	x"065d",	x"06a4",	
												x"069a",	x"067d",	x"069e",	x"0686",	
												x"06a7",	x"0686",	x"06a4",	x"0699",	
												x"0699",	x"068c",	x"06ab",	x"068d",	
												x"06d3",	x"0697",	x"0669",	x"0684",	
												x"1031",	x"101b",	x"066d",	x"0666",	
												x"066c",	x"0649",	x"066c",	x"064d",	
												x"0654",	x"065e",	x"064d",	x"0612",	
												x"0658",	x"064a",	x"0616",	x"0649",	
												x"0618",	x"0662",	x"062d",	x"0628",	
												x"0684",	x"063b",	x"06a6",	x"067b",	
												x"068d",	x"06a8",	x"067f",	x"068e",	
												x"06a5",	x"068f",	x"068d",	x"06a3",	
												x"0642",	x"069d",	x"0664",	x"0652",	
												x"0679",	x"0667",	x"0686",	x"0677",	
												x"0676",	x"06af",	x"068a",	x"066d",	
												x"0692",	x"068d",	x"0678",	x"069a",	
												x"064f",	x"068b",	x"067c",	x"067d",	
												x"0691",	x"0696",	x"0693",	x"067a",	
												x"068b",	x"06a0",	x"069e",	x"0676",	
												x"06a8",	x"0692",	x"06a7",	x"06ae",	
												x"062b",	x"06a0",	x"2031",	x"101b",	
												x"065a",	x"063d",	x"066e",	x"0672",	
												x"0665",	x"0644",	x"0654",	x"0661",	
												x"0629",	x"066f",	x"0645",	x"063f",	
												x"064d",	x"064a",	x"061c",	x"064a",	
												x"062a",	x"062f",	x"0640",	x"0644",	
												x"0672",	x"0648",	x"0687",	x"066b",	
												x"0687",	x"067d",	x"067b",	x"0672",	
												x"0698",	x"0687",	x"0641",	x"0673",	
												x"066b",	x"0637",	x"0689",	x"066c",	
												x"0680",	x"067f",	x"065e",	x"0676",	
												x"0679",	x"0655",	x"068b",	x"0676",	
												x"067e",	x"067d",	x"0669",	x"0685",	
												x"0677",	x"0674",	x"068c",	x"067f",	
												x"0675",	x"068a",	x"068d",	x"0676",	
												x"06aa",	x"066f",	x"068a",	x"0692",	
												x"068f",	x"0673",	x"0637",	x"0677",	
												x"3031",	x"101b",	x"064f",	x"0635",	
												x"0643",	x"0641",	x"063b",	x"0645",	
												x"063d",	x"061a",	x"0650",	x"0624",	
												x"0633",	x"062e",	x"0625",	x"0622",	
												x"061f",	x"061d",	x"063b",	x"061f",	
												x"064c",	x"063e",	x"0671",	x"065a",	
												x"067c",	x"065e",	x"0683",	x"0654",	
												x"0674",	x"066d",	x"0687",	x"066d",	
												x"0650",	x"0669",	x"0662",	x"0636",	
												x"0679",	x"0655",	x"0674",	x"066b",	
												x"0675",	x"067e",	x"0683",	x"0662",	
												x"06a1",	x"067b",	x"069e",	x"0690",	
												x"0684",	x"0692",	x"0696",	x"066c",	
												x"069d",	x"0665",	x"0699",	x"0671",	
												x"069f",	x"0695",	x"06aa",	x"0683",	
												x"06b2",	x"0687",	x"06b4",	x"0686",	
												x"066e",	x"0687",	x"0004",	x"000a",	
												x"d88a",	x"fac7",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"101c",	
												x"0693",	x"0649",	x"067a",	x"065d",	
												x"066f",	x"0649",	x"0664",	x"0655",	
												x"067e",	x"0650",	x"0653",	x"0651",	
												x"0659",	x"0656",	x"065d",	x"064c",	
												x"069a",	x"063c",	x"0671",	x"065f",	
												x"06be",	x"0665",	x"06a4",	x"069a",	
												x"06b3",	x"069e",	x"06e4",	x"069d",	
												x"0696",	x"06ab",	x"069b",	x"0691",	
												x"06c6",	x"0696",	x"06c6",	x"06bb",	
												x"06c7",	x"06b3",	x"06d7",	x"06c1",	
												x"06ce",	x"06ca",	x"06dd",	x"06b5",	
												x"06d0",	x"06be",	x"06a1",	x"06ad",	
												x"06df",	x"06a4",	x"06ca",	x"06b4",	
												x"06de",	x"06ba",	x"06ee",	x"06d0",	
												x"06eb",	x"06ca",	x"06ee",	x"06d3",	
												x"06f1",	x"06ce",	x"069b",	x"06cf",	
												x"5031",	x"101c",	x"06a1",	x"069c",	
												x"06b9",	x"0690",	x"06aa",	x"067d",	
												x"06b8",	x"068a",	x"06ac",	x"0693",	
												x"06a9",	x"067c",	x"06a5",	x"068f",	
												x"06a1",	x"0697",	x"06c8",	x"067a",	
												x"06d6",	x"06b0",	x"06d5",	x"06c8",	
												x"06f6",	x"06d2",	x"0701",	x"06d5",	
												x"06e4",	x"06da",	x"06dd",	x"06bb",	
												x"06d4",	x"06bf",	x"0715",	x"06ab",	
												x"06e2",	x"06ca",	x"06f2",	x"06ba",	
												x"06f8",	x"06e0",	x"06f5",	x"06cb",	
												x"0701",	x"06e1",	x"06fb",	x"06d6",	
												x"06e8",	x"06c8",	x"0725",	x"06c8",	
												x"0726",	x"06d5",	x"0729",	x"06d0",	
												x"071d",	x"06f0",	x"071e",	x"06ec",	
												x"0723",	x"0703",	x"072b",	x"06fc",	
												x"06a3",	x"06f8",	x"6031",	x"101c",	
												x"06d9",	x"06a7",	x"06d0",	x"069d",	
												x"06ae",	x"06a7",	x"06bb",	x"0691",	
												x"06cf",	x"0677",	x"06c8",	x"06a9",	
												x"06d2",	x"0688",	x"068c",	x"0684",	
												x"06f7",	x"0686",	x"06fe",	x"06c1",	
												x"072f",	x"06e0",	x"0732",	x"0712",	
												x"0729",	x"06c2",	x"0721",	x"0713",	
												x"071b",	x"06f9",	x"06e3",	x"06f7",	
												x"0710",	x"06ee",	x"0718",	x"0706",	
												x"0737",	x"0700",	x"0738",	x"070d",	
												x"073e",	x"0707",	x"0732",	x"0710",	
												x"0732",	x"0711",	x"071a",	x"06e7",	
												x"0747",	x"06f2",	x"0743",	x"0715",	
												x"0752",	x"070c",	x"075a",	x"0711",	
												x"075d",	x"0715",	x"0755",	x"0730",	
												x"0741",	x"0723",	x"06e9",	x"0716",	
												x"7031",	x"101c",	x"070a",	x"06d0",	
												x"0716",	x"06f9",	x"0737",	x"06dc",	
												x"0731",	x"0701",	x"0719",	x"06ed",	
												x"0734",	x"070d",	x"070f",	x"06f8",	
												x"0701",	x"06da",	x"0731",	x"06c1",	
												x"074e",	x"071d",	x"076a",	x"0732",	
												x"07a5",	x"0770",	x"078c",	x"0758",	
												x"0799",	x"0777",	x"0784",	x"077a",	
												x"0740",	x"0744",	x"077f",	x"0720",	
												x"0781",	x"075a",	x"079a",	x"0761",	
												x"07a0",	x"0776",	x"07a9",	x"0771",	
												x"07ab",	x"077b",	x"07b8",	x"0781",	
												x"0766",	x"077e",	x"0799",	x"0749",	
												x"07b2",	x"0783",	x"07c1",	x"0799",	
												x"07d7",	x"0792",	x"07cc",	x"0796",	
												x"07da",	x"07b5",	x"07ca",	x"07ad",	
												x"070e",	x"0799",	x"0004",	x"000a",	
												x"227f",	x"344c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"201d",	
												x"0732",	x"072f",	x"071d",	x"073f",	
												x"06fb",	x"0712",	x"0719",	x"0721",	
												x"0707",	x"0717",	x"0717",	x"06e8",	
												x"0719",	x"06fa",	x"0721",	x"06f9",	
												x"0724",	x"0740",	x"0737",	x"074c",	
												x"073c",	x"074d",	x"0748",	x"0760",	
												x"075b",	x"0768",	x"0760",	x"0761",	
												x"0747",	x"075a",	x"070c",	x"0737",	
												x"075a",	x"072d",	x"0754",	x"0774",	
												x"073e",	x"0757",	x"074d",	x"0755",	
												x"0736",	x"0742",	x"074f",	x"0759",	
												x"075a",	x"0758",	x"0732",	x"075f",	
												x"0732",	x"0751",	x"072f",	x"072a",	
												x"074e",	x"0735",	x"074e",	x"0740",	
												x"075e",	x"0744",	x"0765",	x"074a",	
												x"074f",	x"0729",	x"06f0",	x"0758",	
												x"1031",	x"201d",	x"0704",	x"0732",	
												x"06fe",	x"06d9",	x"06f3",	x"0709",	
												x"0709",	x"070d",	x"06e9",	x"06d8",	
												x"0703",	x"06ff",	x"071b",	x"0705",	
												x"06cb",	x"0745",	x"0742",	x"06ec",	
												x"073c",	x"0742",	x"075e",	x"072d",	
												x"0769",	x"0762",	x"074f",	x"074e",	
												x"0765",	x"0760",	x"0731",	x"076b",	
												x"06e5",	x"0745",	x"0703",	x"06f3",	
												x"0755",	x"072c",	x"072a",	x"073b",	
												x"0733",	x"0730",	x"0731",	x"073c",	
												x"0755",	x"0744",	x"073f",	x"0748",	
												x"0734",	x"0752",	x"0743",	x"073f",	
												x"0748",	x"074d",	x"076b",	x"0750",	
												x"076d",	x"075c",	x"0761",	x"0752",	
												x"0773",	x"076b",	x"0760",	x"0769",	
												x"06f3",	x"0752",	x"2031",	x"201d",	
												x"06fe",	x"0717",	x"0705",	x"0721",	
												x"0716",	x"070e",	x"06ed",	x"06fb",	
												x"06e7",	x"06f3",	x"0712",	x"06f2",	
												x"0701",	x"0701",	x"06e5",	x"071b",	
												x"06f2",	x"0700",	x"074f",	x"0736",	
												x"074d",	x"075e",	x"0747",	x"0753",	
												x"0737",	x"0751",	x"0737",	x"0734",	
												x"074f",	x"0732",	x"06fc",	x"0733",	
												x"0749",	x"0700",	x"0713",	x"073b",	
												x"0739",	x"0727",	x"073b",	x"073a",	
												x"074e",	x"073b",	x"0747",	x"073e",	
												x"0745",	x"074d",	x"0704",	x"0742",	
												x"0748",	x"0724",	x"0756",	x"072b",	
												x"0733",	x"072e",	x"073d",	x"073a",	
												x"0768",	x"0731",	x"0769",	x"075d",	
												x"0752",	x"0752",	x"06dd",	x"0744",	
												x"3031",	x"201d",	x"06f9",	x"06f4",	
												x"0707",	x"06d7",	x"0718",	x"06d5",	
												x"06f8",	x"0700",	x"06f5",	x"06eb",	
												x"06df",	x"06eb",	x"070b",	x"06db",	
												x"06ff",	x"0702",	x"0720",	x"06f7",	
												x"0741",	x"070c",	x"0766",	x"071f",	
												x"0761",	x"0753",	x"0756",	x"0757",	
												x"074e",	x"075a",	x"0743",	x"0728",	
												x"06f4",	x"0734",	x"0733",	x"070c",	
												x"073b",	x"072f",	x"075a",	x"073b",	
												x"0771",	x"0762",	x"076e",	x"073f",	
												x"0770",	x"074f",	x"074d",	x"0755",	
												x"0754",	x"073e",	x"0784",	x"073c",	
												x"075c",	x"074b",	x"076b",	x"072b",	
												x"0764",	x"0728",	x"0786",	x"0739",	
												x"0793",	x"074e",	x"0796",	x"075c",	
												x"0724",	x"0758",	x"0004",	x"000a",	
												x"3a02",	x"9d4d",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"201e",	
												x"0730",	x"071a",	x"072e",	x"0742",	
												x"072e",	x"071b",	x"0745",	x"072d",	
												x"070a",	x"0701",	x"073c",	x"0724",	
												x"0741",	x"0700",	x"072c",	x"0720",	
												x"074f",	x"0729",	x"0772",	x"0761",	
												x"0776",	x"0768",	x"07a3",	x"0769",	
												x"0790",	x"075b",	x"0783",	x"0766",	
												x"0773",	x"0781",	x"075a",	x"0764",	
												x"0796",	x"0752",	x"0799",	x"0769",	
												x"07ad",	x"0784",	x"079a",	x"0791",	
												x"07c4",	x"077c",	x"07c4",	x"0796",	
												x"07c2",	x"07aa",	x"0798",	x"079f",	
												x"07c0",	x"0799",	x"07a6",	x"07b8",	
												x"07b9",	x"079e",	x"07a3",	x"078c",	
												x"07c2",	x"0782",	x"07cf",	x"079c",	
												x"07c8",	x"07af",	x"0747",	x"0792",	
												x"5031",	x"201e",	x"076a",	x"0744",	
												x"079d",	x"0748",	x"078b",	x"074b",	
												x"076a",	x"0745",	x"076c",	x"0732",	
												x"0788",	x"074e",	x"077b",	x"0756",	
												x"0792",	x"0755",	x"07c9",	x"0783",	
												x"07d3",	x"0786",	x"07b7",	x"0791",	
												x"07ba",	x"07a7",	x"07d7",	x"07ad",	
												x"07b1",	x"07b6",	x"07bf",	x"07ac",	
												x"0790",	x"0785",	x"07db",	x"0763",	
												x"07e0",	x"0798",	x"07e1",	x"078b",	
												x"07f4",	x"07a0",	x"07dc",	x"0795",	
												x"0802",	x"07c2",	x"07e8",	x"07a5",	
												x"07cc",	x"07b0",	x"07f9",	x"07ab",	
												x"07e4",	x"07c0",	x"07ea",	x"07aa",	
												x"0803",	x"0795",	x"0806",	x"07aa",	
												x"080d",	x"07be",	x"07e3",	x"07c4",	
												x"0765",	x"07a4",	x"6031",	x"201e",	
												x"07a7",	x"0771",	x"0789",	x"0785",	
												x"077a",	x"0760",	x"07a7",	x"0753",	
												x"0774",	x"075c",	x"07c7",	x"0744",	
												x"079e",	x"076d",	x"07ae",	x"077b",	
												x"07fc",	x"0779",	x"0802",	x"07bf",	
												x"07f1",	x"07b2",	x"0807",	x"07bf",	
												x"080a",	x"07be",	x"0800",	x"07eb",	
												x"07e5",	x"07d9",	x"07e7",	x"07d9",	
												x"07f4",	x"07c6",	x"080a",	x"07e6",	
												x"081b",	x"07d7",	x"082a",	x"07f1",	
												x"0823",	x"07df",	x"0833",	x"07f3",	
												x"082f",	x"07e2",	x"0801",	x"07e6",	
												x"0821",	x"07f3",	x"082b",	x"07db",	
												x"0852",	x"07ce",	x"083b",	x"07e6",	
												x"0841",	x"07fc",	x"0842",	x"07fd",	
												x"0838",	x"07fc",	x"07c9",	x"07e8",	
												x"7031",	x"201e",	x"07f7",	x"07b5",	
												x"07d2",	x"07b1",	x"07ef",	x"079d",	
												x"0810",	x"07ac",	x"07f5",	x"07a0",	
												x"081b",	x"0794",	x"0816",	x"079c",	
												x"07f3",	x"07b5",	x"085f",	x"07d7",	
												x"086d",	x"0829",	x"0870",	x"0827",	
												x"087c",	x"0824",	x"088a",	x"082e",	
												x"086c",	x"0856",	x"086a",	x"0843",	
												x"087a",	x"0845",	x"0886",	x"082c",	
												x"08a8",	x"0846",	x"08a0",	x"085b",	
												x"08a2",	x"0858",	x"08a3",	x"0849",	
												x"0887",	x"0867",	x"08d7",	x"0854",	
												x"0881",	x"086f",	x"08a9",	x"087c",	
												x"0896",	x"087f",	x"08b9",	x"0873",	
												x"08b8",	x"0888",	x"08bf",	x"0887",	
												x"08d2",	x"0887",	x"088e",	x"0895",	
												x"06ff",	x"089f",	x"0004",	x"000a",	
												x"92bd",	x"dfbc",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"301f",	
												x"06e6",	x"06f0",	x"0709",	x"06df",	
												x"06ea",	x"06fb",	x"06ef",	x"0727",	
												x"070a",	x"06fa",	x"06fa",	x"06f1",	
												x"06f3",	x"06e2",	x"06c8",	x"06ef",	
												x"06ff",	x"06d9",	x"0730",	x"0723",	
												x"0711",	x"072a",	x"0755",	x"0721",	
												x"075e",	x"073a",	x"075b",	x"0751",	
												x"0711",	x"0743",	x"06de",	x"0711",	
												x"0711",	x"070a",	x"071d",	x"0727",	
												x"06ee",	x"0716",	x"0744",	x"071b",	
												x"0748",	x"0732",	x"0749",	x"0742",	
												x"071d",	x"0715",	x"0718",	x"070f",	
												x"071b",	x"071f",	x"071c",	x"0724",	
												x"070f",	x"070c",	x"070c",	x"070f",	
												x"072f",	x"0701",	x"074f",	x"072d",	
												x"073a",	x"0749",	x"06d0",	x"0713",	
												x"1031",	x"301f",	x"06c6",	x"06f0",	
												x"06cc",	x"06e5",	x"06cf",	x"06c5",	
												x"06d1",	x"06bc",	x"06d1",	x"06bd",	
												x"06d6",	x"06ef",	x"06dd",	x"06c5",	
												x"06b1",	x"06df",	x"0714",	x"06c8",	
												x"073b",	x"071b",	x"0723",	x"0748",	
												x"0719",	x"0737",	x"0711",	x"071c",	
												x"071c",	x"071b",	x"0719",	x"0715",	
												x"06c5",	x"0714",	x"071c",	x"06db",	
												x"0709",	x"0721",	x"0727",	x"0715",	
												x"0739",	x"0736",	x"0720",	x"0748",	
												x"0754",	x"073f",	x"072c",	x"0740",	
												x"0713",	x"072f",	x"070d",	x"070c",	
												x"0739",	x"070d",	x"072f",	x"0743",	
												x"0712",	x"0725",	x"0722",	x"0707",	
												x"0724",	x"0718",	x"0725",	x"0721",	
												x"06dc",	x"073e",	x"2031",	x"301f",	
												x"06d3",	x"06e3",	x"06b7",	x"06d3",	
												x"06bd",	x"06ba",	x"06d6",	x"06cc",	
												x"06cd",	x"06e9",	x"06d5",	x"06c5",	
												x"06e4",	x"06ce",	x"0677",	x"0709",	
												x"0709",	x"06e1",	x"070f",	x"0723",	
												x"071e",	x"071e",	x"0710",	x"0709",	
												x"0728",	x"071f",	x"0723",	x"0723",	
												x"070b",	x"0703",	x"06db",	x"070e",	
												x"0709",	x"0708",	x"070a",	x"0705",	
												x"0703",	x"06fd",	x"071f",	x"0718",	
												x"072b",	x"0719",	x"0746",	x"0725",	
												x"072c",	x"0736",	x"06e6",	x"0720",	
												x"070f",	x"06f1",	x"0739",	x"0721",	
												x"0712",	x"0708",	x"0731",	x"0705",	
												x"0708",	x"0710",	x"071f",	x"0703",	
												x"072e",	x"0709",	x"069f",	x"0722",	
												x"3031",	x"301f",	x"06b0",	x"0696",	
												x"06e5",	x"06a8",	x"06ba",	x"06be",	
												x"070c",	x"06c0",	x"06e2",	x"06c5",	
												x"06d5",	x"06cf",	x"06d5",	x"06cd",	
												x"06de",	x"06c8",	x"06f3",	x"06d6",	
												x"0703",	x"06fd",	x"0727",	x"06f7",	
												x"0724",	x"0710",	x"071f",	x"0705",	
												x"06eb",	x"070d",	x"06f6",	x"06ea",	
												x"06de",	x"070a",	x"06f9",	x"06db",	
												x"06ff",	x"06f1",	x"072c",	x"06f3",	
												x"0733",	x"0727",	x"0726",	x"071e",	
												x"075a",	x"0728",	x"0753",	x"0708",	
												x"0729",	x"0724",	x"0732",	x"0710",	
												x"0718",	x"0717",	x"071a",	x"0702",	
												x"072d",	x"0700",	x"072f",	x"0702",	
												x"0739",	x"0702",	x"072f",	x"06eb",	
												x"06e1",	x"070d",	x"0004",	x"000a",	
												x"246f",	x"c758",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"3020",	
												x"06f7",	x"06b2",	x"06ee",	x"06f2",	
												x"06f0",	x"06cd",	x"0706",	x"06ca",	
												x"06f4",	x"06d9",	x"0700",	x"06ee",	
												x"070f",	x"070e",	x"0707",	x"0709",	
												x"0731",	x"06f8",	x"073f",	x"0736",	
												x"074c",	x"0733",	x"0751",	x"0742",	
												x"0752",	x"073d",	x"075b",	x"0735",	
												x"072c",	x"0739",	x"0708",	x"0717",	
												x"0759",	x"06f9",	x"0754",	x"0740",	
												x"0757",	x"073c",	x"077c",	x"0752",	
												x"0769",	x"0749",	x"0771",	x"074d",	
												x"0774",	x"075c",	x"0743",	x"0757",	
												x"074f",	x"0744",	x"077f",	x"073b",	
												x"075e",	x"0759",	x"076f",	x"0765",	
												x"0779",	x"0751",	x"0783",	x"075c",	
												x"0776",	x"074e",	x"0748",	x"0744",	
												x"5031",	x"3020",	x"074b",	x"0722",	
												x"073b",	x"0727",	x"0748",	x"06f7",	
												x"074c",	x"072b",	x"074f",	x"0720",	
												x"076a",	x"072c",	x"076f",	x"0750",	
												x"075b",	x"0751",	x"077e",	x"0756",	
												x"077a",	x"0788",	x"077b",	x"076a",	
												x"0776",	x"0766",	x"078b",	x"0759",	
												x"077e",	x"0773",	x"0775",	x"0775",	
												x"0750",	x"075b",	x"07a8",	x"0725",	
												x"078d",	x"074d",	x"079b",	x"0769",	
												x"07bd",	x"077f",	x"07b0",	x"0773",	
												x"07c1",	x"0775",	x"07c8",	x"077d",	
												x"07a4",	x"077a",	x"07e1",	x"0759",	
												x"07a6",	x"0785",	x"07b0",	x"0779",	
												x"07a3",	x"0781",	x"07d4",	x"0747",	
												x"07d0",	x"077b",	x"07c1",	x"0793",	
												x"0738",	x"0791",	x"6031",	x"3020",	
												x"0766",	x"070b",	x"0763",	x"073c",	
												x"0762",	x"072e",	x"0757",	x"0744",	
												x"075d",	x"074f",	x"075e",	x"0759",	
												x"0757",	x"0740",	x"0772",	x"074e",	
												x"07bd",	x"0756",	x"07c2",	x"079e",	
												x"07bd",	x"0799",	x"07c7",	x"07b3",	
												x"07b3",	x"07a3",	x"07b8",	x"0777",	
												x"07c7",	x"0785",	x"0790",	x"0789",	
												x"07bc",	x"0785",	x"07e7",	x"078c",	
												x"07ec",	x"078f",	x"07ec",	x"07b7",	
												x"07fd",	x"07b0",	x"0801",	x"07a5",	
												x"07e4",	x"07a8",	x"07c0",	x"07a8",	
												x"07f2",	x"07af",	x"07dc",	x"07d2",	
												x"07e6",	x"07ad",	x"0814",	x"07c1",	
												x"07ff",	x"07ad",	x"0813",	x"07e0",	
												x"0800",	x"07c7",	x"078a",	x"07c8",	
												x"7031",	x"3020",	x"0797",	x"076f",	
												x"07a8",	x"074c",	x"07b1",	x"0760",	
												x"07f5",	x"0780",	x"07b8",	x"078f",	
												x"07d4",	x"077d",	x"07e1",	x"0794",	
												x"07f1",	x"07d3",	x"084a",	x"07cd",	
												x"0842",	x"07e0",	x"082d",	x"0806",	
												x"0823",	x"0800",	x"084b",	x"07f6",	
												x"083b",	x"0827",	x"081c",	x"0807",	
												x"07e4",	x"07f6",	x"083b",	x"07e6",	
												x"0858",	x"0818",	x"0862",	x"0803",	
												x"085c",	x"0839",	x"0868",	x"0818",	
												x"0886",	x"083d",	x"0872",	x"085d",	
												x"082d",	x"0848",	x"086d",	x"082a",	
												x"087d",	x"085b",	x"086a",	x"081d",	
												x"08ba",	x"084e",	x"089e",	x"0854",	
												x"088c",	x"086a",	x"086d",	x"086d",	
												x"06c8",	x"0852",	x"0004",	x"000a",	
												x"754a",	x"05ed",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"0121",	
												x"0669",	x"0665",	x"0655",	x"065c",	
												x"0663",	x"065b",	x"0653",	x"065e",	
												x"0663",	x"064b",	x"065b",	x"0636",	
												x"065c",	x"0662",	x"065d",	x"0659",	
												x"065e",	x"0659",	x"069e",	x"0675",	
												x"0662",	x"0683",	x"0662",	x"067d",	
												x"0672",	x"0658",	x"069d",	x"0686",	
												x"068f",	x"067e",	x"063e",	x"068a",	
												x"0669",	x"0654",	x"0678",	x"0698",	
												x"069c",	x"0675",	x"067f",	x"067d",	
												x"0665",	x"067c",	x"06a5",	x"067b",	
												x"066a",	x"068d",	x"064b",	x"066f",	
												x"0672",	x"065e",	x"06a6",	x"067b",	
												x"0696",	x"068c",	x"06a4",	x"06a1",	
												x"067c",	x"0694",	x"06c2",	x"0682",	
												x"0683",	x"068d",	x"0671",	x"0675",	
												x"102e",	x"0121",	x"063c",	x"0666",	
												x"063e",	x"0655",	x"0640",	x"0632",	
												x"0617",	x"064e",	x"0620",	x"0622",	
												x"0634",	x"062a",	x"063d",	x"0630",	
												x"0623",	x"065b",	x"0656",	x"0650",	
												x"066c",	x"0668",	x"066e",	x"0663",	
												x"0674",	x"066d",	x"0663",	x"068a",	
												x"0678",	x"067f",	x"0678",	x"0683",	
												x"0632",	x"066a",	x"0673",	x"064f",	
												x"0664",	x"067d",	x"064a",	x"065b",	
												x"0678",	x"0669",	x"067f",	x"0683",	
												x"067b",	x"0685",	x"0670",	x"066d",	
												x"0632",	x"0670",	x"0660",	x"0665",	
												x"066e",	x"068b",	x"068a",	x"0684",	
												x"068a",	x"0692",	x"068a",	x"067e",	
												x"068d",	x"06b8",	x"0681",	x"0699",	
												x"0626",	x"0681",	x"202e",	x"0121",	
												x"0629",	x"0623",	x"062a",	x"063c",	
												x"0612",	x"063c",	x"0623",	x"0643",	
												x"0629",	x"063a",	x"0652",	x"064b",	
												x"065d",	x"0657",	x"061f",	x"0663",	
												x"0633",	x"063b",	x"0638",	x"0654",	
												x"0660",	x"0647",	x"064f",	x"0651",	
												x"0674",	x"066e",	x"0682",	x"068a",	
												x"0678",	x"067c",	x"0641",	x"0686",	
												x"0639",	x"0651",	x"0635",	x"065a",	
												x"0654",	x"063d",	x"0654",	x"066a",	
												x"0670",	x"064f",	x"066f",	x"0662",	
												x"0661",	x"065b",	x"063a",	x"064f",	
												x"0658",	x"0656",	x"0645",	x"064e",	
												x"0670",	x"0651",	x"068f",	x"066e",	
												x"065f",	x"067d",	x"068c",	x"0673",	
												x"0679",	x"066a",	x"0615",	x"0660",	
												x"302e",	x"0121",	x"0628",	x"060f",	
												x"061d",	x"0623",	x"061d",	x"0621",	
												x"0602",	x"060f",	x"0627",	x"0601",	
												x"0639",	x"0630",	x"062b",	x"0636",	
												x"061a",	x"0634",	x"064c",	x"063b",	
												x"0660",	x"0662",	x"065c",	x"064a",	
												x"0649",	x"0661",	x"0644",	x"063a",	
												x"0667",	x"0653",	x"064a",	x"0651",	
												x"0621",	x"0654",	x"063f",	x"063a",	
												x"064e",	x"0651",	x"0643",	x"0642",	
												x"0669",	x"0665",	x"0681",	x"0661",	
												x"0661",	x"0677",	x"0677",	x"065e",	
												x"0643",	x"0652",	x"0666",	x"064e",	
												x"0687",	x"0659",	x"0676",	x"065d",	
												x"0672",	x"0672",	x"0686",	x"0668",	
												x"0687",	x"066c",	x"0675",	x"065b",	
												x"0626",	x"0661",	x"0004",	x"000a",	
												x"cd8c",	x"b865",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"0122",	
												x"063a",	x"0613",	x"0653",	x"0636",	
												x"061a",	x"0619",	x"062e",	x"062a",	
												x"0638",	x"063c",	x"0661",	x"063b",	
												x"0656",	x"0654",	x"0654",	x"0642",	
												x"0654",	x"0659",	x"067b",	x"065a",	
												x"065e",	x"0651",	x"0666",	x"0676",	
												x"067a",	x"0668",	x"066f",	x"0663",	
												x"0677",	x"0680",	x"0652",	x"067b",	
												x"066f",	x"065d",	x"0682",	x"0677",	
												x"068f",	x"067b",	x"068c",	x"0699",	
												x"0696",	x"0689",	x"069b",	x"06a4",	
												x"065f",	x"0689",	x"067c",	x"0680",	
												x"067a",	x"068c",	x"06a2",	x"0689",	
												x"06a7",	x"06a3",	x"069d",	x"06c1",	
												x"06ad",	x"0691",	x"06ba",	x"06a6",	
												x"06a4",	x"06a3",	x"066e",	x"069b",	
												x"502e",	x"0122",	x"0689",	x"0659",	
												x"0655",	x"0673",	x"064f",	x"0647",	
												x"066e",	x"0640",	x"0676",	x"0641",	
												x"0668",	x"0668",	x"0694",	x"0667",	
												x"066b",	x"0681",	x"069a",	x"0682",	
												x"069f",	x"068c",	x"0693",	x"0691",	
												x"06ac",	x"069c",	x"069b",	x"06a1",	
												x"069b",	x"06a7",	x"06a3",	x"0699",	
												x"0680",	x"0692",	x"0688",	x"066b",	
												x"06af",	x"069a",	x"06a2",	x"068f",	
												x"06ab",	x"069d",	x"06b5",	x"06b2",	
												x"06ad",	x"068f",	x"06b1",	x"06a7",	
												x"06a3",	x"06a3",	x"06ca",	x"0696",	
												x"06d5",	x"06b3",	x"06e2",	x"06bd",	
												x"06e4",	x"06ad",	x"06d5",	x"06b9",	
												x"06da",	x"06b0",	x"06c8",	x"06bc",	
												x"0671",	x"06b1",	x"602e",	x"0122",	
												x"0686",	x"065b",	x"0689",	x"066c",	
												x"0653",	x"0673",	x"0667",	x"0663",	
												x"06a2",	x"066b",	x"067b",	x"06ab",	
												x"067d",	x"0668",	x"067a",	x"068f",	
												x"068f",	x"066f",	x"06c4",	x"067e",	
												x"069e",	x"06a2",	x"06cf",	x"06a5",	
												x"06d2",	x"06d2",	x"06fc",	x"06cc",	
												x"06c9",	x"06cb",	x"06b2",	x"06d3",	
												x"06c7",	x"06a6",	x"06d4",	x"06c1",	
												x"06df",	x"06b3",	x"06e2",	x"06d9",	
												x"06ec",	x"06dd",	x"06e4",	x"06e0",	
												x"06f1",	x"06d3",	x"06c7",	x"06c6",	
												x"0709",	x"06d6",	x"0700",	x"0700",	
												x"0709",	x"06e6",	x"0702",	x"06f3",	
												x"070a",	x"06db",	x"0713",	x"06f4",	
												x"0702",	x"06eb",	x"069c",	x"06ec",	
												x"702e",	x"0122",	x"0696",	x"065a",	
												x"0699",	x"0688",	x"068e",	x"0673",	
												x"06a1",	x"0678",	x"06b4",	x"067d",	
												x"06c2",	x"069e",	x"0694",	x"06c8",	
												x"06c2",	x"0686",	x"06c2",	x"06a3",	
												x"071c",	x"0706",	x"06f9",	x"06f8",	
												x"071a",	x"06d6",	x"073b",	x"06f9",	
												x"0741",	x"0714",	x"0723",	x"06fa",	
												x"06e7",	x"071f",	x"074b",	x"06ea",	
												x"0722",	x"071c",	x"073c",	x"0724",	
												x"0754",	x"0737",	x"0757",	x"0747",	
												x"073e",	x"0746",	x"0743",	x"072d",	
												x"0729",	x"0730",	x"074e",	x"0738",	
												x"076a",	x"074b",	x"074a",	x"075c",	
												x"0777",	x"075a",	x"0776",	x"0764",	
												x"0780",	x"075b",	x"0769",	x"0756",	
												x"071b",	x"0754",	x"0004",	x"000a",	
												x"fcdd",	x"deab",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"1123",	
												x"0729",	x"0711",	x"0733",	x"0710",	
												x"0700",	x"0725",	x"06fa",	x"071b",	
												x"0728",	x"0712",	x"076a",	x"0720",	
												x"0762",	x"074d",	x"0726",	x"0750",	
												x"075f",	x"0728",	x"0789",	x"0772",	
												x"077a",	x"0776",	x"076e",	x"077a",	
												x"0734",	x"0750",	x"0745",	x"0750",	
												x"074b",	x"0750",	x"072f",	x"0774",	
												x"0748",	x"074f",	x"075e",	x"0755",	
												x"0742",	x"0755",	x"0742",	x"074c",	
												x"0740",	x"0747",	x"075e",	x"074d",	
												x"0750",	x"075b",	x"070d",	x"0748",	
												x"0767",	x"076b",	x"075e",	x"0772",	
												x"0762",	x"075c",	x"0769",	x"0767",	
												x"0750",	x"075e",	x"0787",	x"0771",	
												x"075d",	x"074c",	x"06ec",	x"0741",	
												x"102e",	x"1123",	x"06f8",	x"06e6",	
												x"0722",	x"073b",	x"0715",	x"0726",	
												x"0704",	x"071a",	x"0700",	x"070d",	
												x"0710",	x"06fe",	x"073b",	x"0719",	
												x"0713",	x"0743",	x"0749",	x"0723",	
												x"074e",	x"074c",	x"0752",	x"073e",	
												x"0737",	x"0744",	x"072c",	x"0739",	
												x"074c",	x"073e",	x"073a",	x"0743",	
												x"0726",	x"073a",	x"0742",	x"0728",	
												x"0750",	x"076d",	x"0758",	x"0743",	
												x"071e",	x"0750",	x"0722",	x"0735",	
												x"073f",	x"071f",	x"0756",	x"0738",	
												x"071f",	x"0767",	x"0753",	x"0749",	
												x"0768",	x"075a",	x"0762",	x"0752",	
												x"0742",	x"075a",	x"0737",	x"075d",	
												x"0744",	x"074d",	x"0758",	x"0740",	
												x"070c",	x"0748",	x"202e",	x"1123",	
												x"06fb",	x"06f3",	x"0702",	x"06f8",	
												x"06d4",	x"0706",	x"0718",	x"06ee",	
												x"06fb",	x"071d",	x"06e9",	x"0726",	
												x"06f7",	x"070e",	x"06e4",	x"0724",	
												x"0732",	x"070a",	x"072c",	x"075a",	
												x"0726",	x"0743",	x"0719",	x"072e",	
												x"0718",	x"072b",	x"0715",	x"072f",	
												x"071d",	x"0725",	x"06f9",	x"073b",	
												x"072d",	x"0713",	x"0724",	x"072b",	
												x"071d",	x"0727",	x"0707",	x"0728",	
												x"0724",	x"070b",	x"071f",	x"071f",	
												x"0730",	x"071b",	x"071a",	x"073f",	
												x"0734",	x"0736",	x"0735",	x"072f",	
												x"072d",	x"073b",	x"0736",	x"0739",	
												x"0734",	x"0726",	x"0731",	x"072d",	
												x"0725",	x"072b",	x"06c6",	x"0710",	
												x"302e",	x"1123",	x"06cf",	x"06b8",	
												x"06e4",	x"06b7",	x"06d5",	x"06d2",	
												x"06ec",	x"06c9",	x"06e1",	x"06ed",	
												x"06b8",	x"06ef",	x"0719",	x"06ca",	
												x"06e6",	x"0707",	x"071e",	x"06f4",	
												x"071c",	x"0719",	x"072b",	x"070d",	
												x"06f3",	x"070d",	x"0727",	x"0718",	
												x"0730",	x"071f",	x"0722",	x"0731",	
												x"06fb",	x"0711",	x"0729",	x"06ff",	
												x"0727",	x"0713",	x"0721",	x"0718",	
												x"071d",	x"0718",	x"071d",	x"0719",	
												x"0731",	x"0702",	x"074c",	x"0713",	
												x"06fa",	x"072a",	x"0728",	x"0732",	
												x"0743",	x"0733",	x"0739",	x"0719",	
												x"073f",	x"072b",	x"0753",	x"0734",	
												x"075c",	x"0730",	x"0755",	x"0723",	
												x"06e8",	x"072f",	x"0004",	x"000a",	
												x"34b0",	x"5f05",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"1124",	
												x"06f8",	x"06d3",	x"0702",	x"06ec",	
												x"06ed",	x"06ef",	x"0706",	x"06fc",	
												x"0704",	x"06ed",	x"0700",	x"0702",	
												x"0710",	x"0715",	x"0704",	x"071c",	
												x"0716",	x"071d",	x"0737",	x"071a",	
												x"0740",	x"073e",	x"0745",	x"0732",	
												x"073a",	x"073e",	x"0742",	x"073e",	
												x"074b",	x"0749",	x"073d",	x"0750",	
												x"0753",	x"0751",	x"0754",	x"0780",	
												x"077f",	x"0747",	x"075d",	x"0766",	
												x"075b",	x"076c",	x"0753",	x"0751",	
												x"074f",	x"0760",	x"0751",	x"0748",	
												x"076b",	x"075d",	x"078b",	x"0761",	
												x"077a",	x"0771",	x"078c",	x"076b",	
												x"078e",	x"0775",	x"07a6",	x"0776",	
												x"0771",	x"0776",	x"073d",	x"074f",	
												x"502e",	x"1124",	x"072b",	x"071c",	
												x"0742",	x"0700",	x"0750",	x"0711",	
												x"0747",	x"0709",	x"0747",	x"0721",	
												x"073e",	x"073b",	x"074c",	x"072b",	
												x"074f",	x"074b",	x"077b",	x"074c",	
												x"0783",	x"0760",	x"076b",	x"0750",	
												x"0771",	x"0765",	x"077a",	x"0774",	
												x"076d",	x"076d",	x"077e",	x"0764",	
												x"0769",	x"076f",	x"077b",	x"075c",	
												x"078c",	x"077e",	x"077a",	x"076b",	
												x"0785",	x"0763",	x"079e",	x"076a",	
												x"07a7",	x"077d",	x"07a3",	x"0778",	
												x"0794",	x"077d",	x"07b8",	x"077a",	
												x"07ae",	x"078a",	x"07bd",	x"0781",	
												x"07c3",	x"078e",	x"07b6",	x"078c",	
												x"07d3",	x"078c",	x"07ad",	x"079e",	
												x"073c",	x"077e",	x"602e",	x"1124",	
												x"072e",	x"0719",	x"074d",	x"06fa",	
												x"0756",	x"0728",	x"075f",	x"0732",	
												x"0747",	x"0735",	x"0760",	x"070a",	
												x"075b",	x"0748",	x"0774",	x"0743",	
												x"077c",	x"0764",	x"078f",	x"0756",	
												x"07b4",	x"0770",	x"07b4",	x"077f",	
												x"07ab",	x"0775",	x"0793",	x"077b",	
												x"0794",	x"077a",	x"079e",	x"0784",	
												x"079e",	x"078d",	x"07b8",	x"07a8",	
												x"07b6",	x"07a0",	x"07af",	x"07c3",	
												x"07bf",	x"07c0",	x"07cc",	x"07ac",	
												x"07ac",	x"07a9",	x"07c6",	x"079f",	
												x"07eb",	x"07bd",	x"07e4",	x"07dd",	
												x"07bc",	x"07bc",	x"07f1",	x"07a4",	
												x"07f7",	x"07cd",	x"07e4",	x"07c1",	
												x"07e2",	x"07bd",	x"076d",	x"0791",	
												x"702e",	x"1124",	x"078b",	x"0761",	
												x"077b",	x"0768",	x"078f",	x"0744",	
												x"0789",	x"0770",	x"0780",	x"0743",	
												x"07af",	x"076d",	x"079e",	x"07a9",	
												x"07ab",	x"0797",	x"07b7",	x"0796",	
												x"07ea",	x"07b4",	x"07f1",	x"07c4",	
												x"0803",	x"07e6",	x"07f1",	x"07cb",	
												x"080d",	x"07f3",	x"07ed",	x"07e9",	
												x"07e8",	x"07ec",	x"07f9",	x"07e6",	
												x"07ef",	x"07eb",	x"083e",	x"07e6",	
												x"0848",	x"07f4",	x"0821",	x"07fd",	
												x"081d",	x"080e",	x"082c",	x"081a",	
												x"07e9",	x"0835",	x"0864",	x"0800",	
												x"0869",	x"0826",	x"083f",	x"0830",	
												x"0867",	x"0843",	x"0891",	x"082c",	
												x"0851",	x"0837",	x"0842",	x"0844",	
												x"06ed",	x"0821",	x"0004",	x"000a",	
												x"69ee",	x"8765",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"2125",	
												x"06c9",	x"06db",	x"06b3",	x"06bf",	
												x"0694",	x"06a6",	x"06b6",	x"06a5",	
												x"06d4",	x"06c4",	x"06fa",	x"06e1",	
												x"06d8",	x"0728",	x"06e1",	x"06e8",	
												x"06f7",	x"06d6",	x"0710",	x"06fd",	
												x"070c",	x"06eb",	x"0717",	x"0728",	
												x"0706",	x"0714",	x"06f0",	x"06ff",	
												x"06f8",	x"06fa",	x"06d7",	x"06f8",	
												x"06f1",	x"070d",	x"06ee",	x"070b",	
												x"06f5",	x"0702",	x"06f3",	x"0715",	
												x"06f1",	x"06f4",	x"06f9",	x"0700",	
												x"06fa",	x"06ff",	x"06f5",	x"06ec",	
												x"0722",	x"06f2",	x"0705",	x"0715",	
												x"071e",	x"0700",	x"072c",	x"06f8",	
												x"0708",	x"070f",	x"06fc",	x"06f5",	
												x"0701",	x"06e6",	x"06a4",	x"06f1",	
												x"102e",	x"2125",	x"0690",	x"069d",	
												x"06b9",	x"068c",	x"06a3",	x"06c0",	
												x"0692",	x"06a5",	x"06b2",	x"0683",	
												x"06d5",	x"06ce",	x"06e1",	x"06be",	
												x"06b4",	x"06b3",	x"06e6",	x"06d3",	
												x"06ec",	x"06e1",	x"06df",	x"06ed",	
												x"06de",	x"06d3",	x"06d9",	x"06de",	
												x"06d9",	x"06e0",	x"06ce",	x"06eb",	
												x"06c1",	x"06f4",	x"06e8",	x"06c5",	
												x"06df",	x"06e5",	x"06e3",	x"06f1",	
												x"06e5",	x"0706",	x"06ee",	x"06fa",	
												x"06eb",	x"0717",	x"06ed",	x"06d5",	
												x"06e2",	x"06fe",	x"070c",	x"06fc",	
												x"0707",	x"0738",	x"0709",	x"0701",	
												x"06dc",	x"0717",	x"0715",	x"06e1",	
												x"0712",	x"0704",	x"06f8",	x"070d",	
												x"06a8",	x"06e5",	x"202e",	x"2125",	
												x"0691",	x"069e",	x"06a6",	x"0695",	
												x"0681",	x"06a3",	x"06ae",	x"06a1",	
												x"06a4",	x"06d1",	x"06aa",	x"06be",	
												x"06a0",	x"069c",	x"0689",	x"06b3",	
												x"06c1",	x"069a",	x"06c0",	x"06ea",	
												x"06d9",	x"06ce",	x"06d8",	x"06ef",	
												x"06d6",	x"06d6",	x"06df",	x"06da",	
												x"06e2",	x"06e0",	x"06ac",	x"06c6",	
												x"06ca",	x"06bd",	x"06ea",	x"06dd",	
												x"06de",	x"06c7",	x"06da",	x"06ef",	
												x"06db",	x"06cd",	x"06e6",	x"06da",	
												x"06dd",	x"06e9",	x"06c6",	x"06c5",	
												x"06e4",	x"06cd",	x"06f8",	x"06de",	
												x"06ee",	x"06e9",	x"06fc",	x"06f5",	
												x"06e5",	x"06ce",	x"06e3",	x"06cf",	
												x"06c5",	x"06cd",	x"0662",	x"06cc",	
												x"302e",	x"2125",	x"0675",	x"0686",	
												x"0680",	x"0667",	x"068f",	x"066a",	
												x"06ac",	x"0695",	x"06ae",	x"068f",	
												x"069a",	x"0699",	x"06aa",	x"06a4",	
												x"0693",	x"06a8",	x"06c5",	x"0696",	
												x"06e9",	x"06bf",	x"06c4",	x"06e7",	
												x"06cf",	x"06c1",	x"06c7",	x"06b3",	
												x"06cd",	x"06d4",	x"06cc",	x"06c9",	
												x"0692",	x"06c0",	x"06cf",	x"06a7",	
												x"06dc",	x"06d8",	x"06d2",	x"06e2",	
												x"06c5",	x"06e3",	x"06ce",	x"06c5",	
												x"06e1",	x"06d3",	x"06e7",	x"06d4",	
												x"06bb",	x"06c0",	x"06f5",	x"06db",	
												x"06f4",	x"06de",	x"06e8",	x"06e6",	
												x"0704",	x"06e1",	x"06ef",	x"06e5",	
												x"06f6",	x"06de",	x"06f0",	x"06d9",	
												x"067d",	x"06d3",	x"0004",	x"000a",	
												x"0a63",	x"7415",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"2126",	
												x"0688",	x"066d",	x"06bb",	x"06a9",	
												x"06a5",	x"06b2",	x"06ab",	x"06a5",	
												x"06ca",	x"06b3",	x"06c2",	x"06ab",	
												x"06e0",	x"06a6",	x"069e",	x"06d1",	
												x"06df",	x"06ae",	x"06e6",	x"06ca",	
												x"06cb",	x"0701",	x"0715",	x"06e8",	
												x"06fc",	x"070b",	x"06fe",	x"06fa",	
												x"06e7",	x"0707",	x"06d1",	x"06f1",	
												x"06f7",	x"06da",	x"071a",	x"071d",	
												x"0704",	x"071a",	x"06fe",	x"0707",	
												x"0707",	x"072e",	x"06f9",	x"0701",	
												x"0705",	x"0701",	x"06fc",	x"06fc",	
												x"071a",	x"0704",	x"071d",	x"0725",	
												x"0734",	x"0709",	x"0724",	x"0732",	
												x"0726",	x"0720",	x"0730",	x"0728",	
												x"072b",	x"071f",	x"06a9",	x"0719",	
												x"502e",	x"2126",	x"06d8",	x"06af",	
												x"06df",	x"06c7",	x"06da",	x"06d9",	
												x"06f7",	x"06cb",	x"0701",	x"06eb",	
												x"06f9",	x"06e9",	x"0708",	x"06f7",	
												x"06e8",	x"0707",	x"0701",	x"06ea",	
												x"072e",	x"06f7",	x"0715",	x"070f",	
												x"071e",	x"073f",	x"070f",	x"0717",	
												x"071a",	x"0718",	x"0715",	x"06fe",	
												x"06f9",	x"0703",	x"0717",	x"06f2",	
												x"071b",	x"0730",	x"071f",	x"070f",	
												x"073b",	x"0712",	x"073d",	x"0702",	
												x"0743",	x"071c",	x"0742",	x"0725",	
												x"073e",	x"0739",	x"0747",	x"0729",	
												x"0740",	x"0732",	x"0750",	x"072c",	
												x"0755",	x"072e",	x"0749",	x"073a",	
												x"0759",	x"073f",	x"076b",	x"072d",	
												x"06d2",	x"073a",	x"602e",	x"2126",	
												x"06d4",	x"06a0",	x"071c",	x"06d6",	
												x"06f0",	x"06f5",	x"06f0",	x"06f0",	
												x"06f5",	x"06d6",	x"071d",	x"06f6",	
												x"06f6",	x"06fc",	x"06d8",	x"06f3",	
												x"072d",	x"06f9",	x"072d",	x"0723",	
												x"0736",	x"0729",	x"0739",	x"0729",	
												x"0762",	x"0722",	x"0755",	x"074d",	
												x"0739",	x"0742",	x"0725",	x"0723",	
												x"074e",	x"071c",	x"0768",	x"0752",	
												x"072d",	x"0742",	x"0763",	x"073d",	
												x"0762",	x"0754",	x"0774",	x"075a",	
												x"0766",	x"0748",	x"0759",	x"0737",	
												x"0789",	x"0749",	x"0790",	x"075f",	
												x"0778",	x"0761",	x"0796",	x"075e",	
												x"079c",	x"0756",	x"0794",	x"0775",	
												x"0791",	x"075c",	x"072c",	x"0749",	
												x"702e",	x"2126",	x"0705",	x"06ef",	
												x"0714",	x"06c0",	x"0724",	x"06f6",	
												x"076f",	x"0722",	x"070a",	x"0718",	
												x"0731",	x"0706",	x"0763",	x"0720",	
												x"0758",	x"071a",	x"0778",	x"0752",	
												x"0791",	x"0764",	x"0790",	x"077c",	
												x"07a2",	x"079f",	x"0790",	x"076c",	
												x"07e1",	x"078c",	x"078e",	x"0778",	
												x"0772",	x"076c",	x"0796",	x"0779",	
												x"07bd",	x"07b2",	x"07c4",	x"07ab",	
												x"07eb",	x"07ba",	x"07c4",	x"07b7",	
												x"07c1",	x"07a9",	x"07d0",	x"07a1",	
												x"07d6",	x"07a3",	x"07ec",	x"07bf",	
												x"07e9",	x"07e2",	x"07f4",	x"07ea",	
												x"0817",	x"07f1",	x"0819",	x"07eb",	
												x"0817",	x"07e6",	x"0808",	x"07dc",	
												x"06de",	x"07ca",	x"0004",	x"000a",	
												x"3ce5",	x"9d2b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"3127",	
												x"070c",	x"06e7",	x"070b",	x"0717",	
												x"06ef",	x"070a",	x"070b",	x"06ef",	
												x"0707",	x"0713",	x"070d",	x"070e",	
												x"0718",	x"071d",	x"0700",	x"0721",	
												x"072d",	x"0729",	x"0729",	x"072c",	
												x"072a",	x"0730",	x"075f",	x"0777",	
												x"075e",	x"073f",	x"0730",	x"0751",	
												x"0719",	x"073c",	x"06f8",	x"070c",	
												x"0722",	x"06f8",	x"0758",	x"073a",	
												x"0753",	x"0754",	x"073d",	x"0759",	
												x"0741",	x"072f",	x"075f",	x"0750",	
												x"073b",	x"0770",	x"06d4",	x"0716",	
												x"072c",	x"0710",	x"0750",	x"0740",	
												x"074f",	x"0730",	x"0777",	x"0761",	
												x"0752",	x"0764",	x"0760",	x"0744",	
												x"072b",	x"0726",	x"06d7",	x"0721",	
												x"102e",	x"3127",	x"06dd",	x"06e7",	
												x"06dc",	x"06f6",	x"06cb",	x"06e1",	
												x"06e9",	x"06f7",	x"06d2",	x"06f0",	
												x"0701",	x"0701",	x"0716",	x"0712",	
												x"06d3",	x"0704",	x"074c",	x"0713",	
												x"0742",	x"073b",	x"073b",	x"0749",	
												x"074b",	x"0759",	x"072d",	x"074e",	
												x"0736",	x"075b",	x"0717",	x"0737",	
												x"06c3",	x"0723",	x"0717",	x"06e3",	
												x"0709",	x"0740",	x"0735",	x"072d",	
												x"072b",	x"0754",	x"071f",	x"0729",	
												x"0714",	x"072d",	x"0727",	x"0721",	
												x"071a",	x"0732",	x"0730",	x"072c",	
												x"0732",	x"072e",	x"072f",	x"0747",	
												x"0750",	x"0740",	x"0745",	x"0745",	
												x"0740",	x"0739",	x"072b",	x"0740",	
												x"06eb",	x"0733",	x"202e",	x"3127",	
												x"06c4",	x"06e5",	x"06c4",	x"06fd",	
												x"06c0",	x"06ff",	x"06e6",	x"06d9",	
												x"06d3",	x"06f5",	x"06f9",	x"06fc",	
												x"06b4",	x"0717",	x"06a9",	x"0708",	
												x"0710",	x"06d2",	x"0710",	x"0736",	
												x"0703",	x"0729",	x"0712",	x"0713",	
												x"0715",	x"071c",	x"0724",	x"0729",	
												x"06fe",	x"06ef",	x"06b6",	x"070c",	
												x"070a",	x"0707",	x"070d",	x"0721",	
												x"0715",	x"071a",	x"0719",	x"06f7",	
												x"071a",	x"070c",	x"0738",	x"071a",	
												x"071f",	x"0712",	x"06be",	x"06f2",	
												x"071c",	x"06e5",	x"071e",	x"072b",	
												x"0715",	x"0739",	x"0713",	x"0727",	
												x"0748",	x"0722",	x"0742",	x"0728",	
												x"070e",	x"0707",	x"06bf",	x"06df",	
												x"302e",	x"3127",	x"06d3",	x"06ac",	
												x"06e5",	x"06ba",	x"06cc",	x"06cf",	
												x"06bd",	x"06c5",	x"06da",	x"06c8",	
												x"06df",	x"06c3",	x"06e3",	x"06c6",	
												x"06e3",	x"06e7",	x"06d9",	x"06d1",	
												x"070e",	x"06dc",	x"0708",	x"06f6",	
												x"0710",	x"06ef",	x"0705",	x"06fe",	
												x"070c",	x"06fa",	x"0709",	x"06fd",	
												x"06ce",	x"0704",	x"06f0",	x"06e5",	
												x"0705",	x"0706",	x"071a",	x"0712",	
												x"0708",	x"071c",	x"071f",	x"0721",	
												x"071c",	x"070d",	x"06fe",	x"070a",	
												x"070a",	x"0702",	x"0702",	x"070e",	
												x"0720",	x"0725",	x"0725",	x"0708",	
												x"0722",	x"0706",	x"0734",	x"0726",	
												x"073d",	x"071e",	x"0729",	x"0719",	
												x"06bc",	x"070e",	x"0004",	x"000a",	
												x"274e",	x"d344",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"3128",	
												x"06d4",	x"06b7",	x"06d1",	x"06bc",	
												x"06cf",	x"06ca",	x"06d6",	x"06d2",	
												x"0700",	x"06c6",	x"0704",	x"06e0",	
												x"06ff",	x"0708",	x"070a",	x"0711",	
												x"0718",	x"06fc",	x"0727",	x"0729",	
												x"0726",	x"071a",	x"0739",	x"0737",	
												x"072d",	x"070f",	x"0726",	x"072d",	
												x"0712",	x"0718",	x"072a",	x"06f1",	
												x"072c",	x"0706",	x"0730",	x"0732",	
												x"0733",	x"072d",	x"0759",	x"0756",	
												x"0748",	x"0746",	x"073c",	x"0751",	
												x"0734",	x"0729",	x"0734",	x"072b",	
												x"0740",	x"073d",	x"075f",	x"0745",	
												x"075e",	x"0754",	x"078a",	x"0779",	
												x"075d",	x"0758",	x"0756",	x"075d",	
												x"0763",	x"0743",	x"0708",	x"0756",	
												x"502e",	x"3128",	x"0701",	x"06d1",	
												x"0713",	x"0700",	x"0716",	x"0703",	
												x"06ff",	x"070d",	x"0734",	x"0707",	
												x"0753",	x"0723",	x"075a",	x"0764",	
												x"0705",	x"0753",	x"0755",	x"0726",	
												x"0758",	x"0756",	x"0760",	x"074f",	
												x"0767",	x"076c",	x"0775",	x"0744",	
												x"074d",	x"0764",	x"0739",	x"074f",	
												x"071f",	x"0734",	x"0772",	x"0726",	
												x"077b",	x"0763",	x"0770",	x"0754",	
												x"078a",	x"077a",	x"0767",	x"076c",	
												x"077e",	x"0765",	x"0766",	x"0760",	
												x"0760",	x"0732",	x"07b6",	x"0750",	
												x"07af",	x"0773",	x"07b1",	x"076a",	
												x"07b8",	x"0778",	x"078f",	x"078f",	
												x"07b4",	x"0763",	x"076e",	x"0775",	
												x"0722",	x"0732",	x"602e",	x"3128",	
												x"0745",	x"0705",	x"0737",	x"06df",	
												x"0736",	x"0730",	x"0738",	x"0714",	
												x"0766",	x"070c",	x"074a",	x"074f",	
												x"0740",	x"0738",	x"072d",	x"072d",	
												x"0783",	x"0722",	x"0783",	x"077c",	
												x"078f",	x"076c",	x"0794",	x"0772",	
												x"0790",	x"077c",	x"0797",	x"0754",	
												x"0787",	x"0762",	x"0785",	x"0760",	
												x"0786",	x"0760",	x"0791",	x"0788",	
												x"0796",	x"0779",	x"07c0",	x"0787",	
												x"079d",	x"077c",	x"07c0",	x"0790",	
												x"07ab",	x"0792",	x"0788",	x"07a0",	
												x"07e7",	x"078b",	x"07e8",	x"07be",	
												x"07dd",	x"07b5",	x"07cf",	x"07bb",	
												x"07d9",	x"079d",	x"07c3",	x"0789",	
												x"07c5",	x"077d",	x"074d",	x"0781",	
												x"702e",	x"3128",	x"075c",	x"0755",	
												x"0772",	x"0748",	x"0755",	x"0756",	
												x"0788",	x"074b",	x"0787",	x"0733",	
												x"07b3",	x"073d",	x"078c",	x"079e",	
												x"078d",	x"0777",	x"07ca",	x"0785",	
												x"080d",	x"07ad",	x"07ca",	x"07ce",	
												x"07f5",	x"07b0",	x"07e6",	x"07b2",	
												x"07e4",	x"07e1",	x"07c9",	x"07dc",	
												x"07ec",	x"07ae",	x"07f5",	x"07db",	
												x"0808",	x"0801",	x"07fd",	x"07fa",	
												x"0844",	x"07fa",	x"0813",	x"07e1",	
												x"080a",	x"080b",	x"07fe",	x"07da",	
												x"080e",	x"07f6",	x"080c",	x"080e",	
												x"0834",	x"080e",	x"0828",	x"0826",	
												x"0868",	x"0822",	x"0856",	x"0814",	
												x"0844",	x"0838",	x"082f",	x"07fe",	
												x"065e",	x"0800",	x"0004",	x"000a",	
												x"5d5b",	x"fb3b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"0129",	
												x"067b",	x"0668",	x"0686",	x"0678",	
												x"0667",	x"067a",	x"066c",	x"0643",	
												x"0656",	x"065a",	x"0644",	x"063f",	
												x"0641",	x"062e",	x"0644",	x"0661",	
												x"0660",	x"0654",	x"0685",	x"0665",	
												x"069f",	x"066e",	x"0695",	x"06ad",	
												x"0689",	x"068c",	x"0691",	x"068e",	
												x"0688",	x"0695",	x"063d",	x"069c",	
												x"0688",	x"0670",	x"0683",	x"0685",	
												x"0697",	x"0683",	x"068b",	x"069d",	
												x"0691",	x"067f",	x"0693",	x"0695",	
												x"0699",	x"069a",	x"063c",	x"0692",	
												x"0692",	x"0678",	x"0695",	x"06b1",	
												x"06a5",	x"06b2",	x"068a",	x"06ad",	
												x"0694",	x"066e",	x"06aa",	x"069c",	
												x"06a8",	x"06ac",	x"0667",	x"0695",	
												x"102f",	x"0129",	x"0626",	x"0654",	
												x"0661",	x"0646",	x"0651",	x"063d",	
												x"0633",	x"0640",	x"0637",	x"063a",	
												x"063a",	x"0623",	x"063d",	x"0626",	
												x"0620",	x"063a",	x"0653",	x"064e",	
												x"068e",	x"0666",	x"0688",	x"068a",	
												x"066a",	x"0678",	x"0689",	x"068f",	
												x"0682",	x"0690",	x"0669",	x"0673",	
												x"064a",	x"066e",	x"0684",	x"064d",	
												x"0675",	x"067d",	x"0678",	x"067d",	
												x"0696",	x"0696",	x"068d",	x"06a6",	
												x"067a",	x"0685",	x"068c",	x"068b",	
												x"063a",	x"0696",	x"067a",	x"067e",	
												x"0688",	x"068b",	x"0689",	x"069a",	
												x"067b",	x"0688",	x"068b",	x"0668",	
												x"069f",	x"06a2",	x"068d",	x"06a4",	
												x"063e",	x"06ac",	x"202f",	x"0129",	
												x"0642",	x"062f",	x"066a",	x"0640",	
												x"064a",	x"0659",	x"0659",	x"064f",	
												x"0620",	x"0655",	x"062d",	x"061e",	
												x"061e",	x"0631",	x"05f4",	x"0642",	
												x"0658",	x"063f",	x"0657",	x"067b",	
												x"0666",	x"0665",	x"066a",	x"0671",	
												x"0665",	x"066e",	x"0671",	x"067c",	
												x"0689",	x"0673",	x"063a",	x"066c",	
												x"0665",	x"0654",	x"0676",	x"0660",	
												x"067a",	x"0668",	x"065a",	x"06a1",	
												x"066d",	x"0667",	x"065b",	x"065b",	
												x"0662",	x"065e",	x"065d",	x"0661",	
												x"0675",	x"066e",	x"066e",	x"0667",	
												x"066f",	x"0668",	x"068f",	x"0678",	
												x"0679",	x"067f",	x"0698",	x"0680",	
												x"0697",	x"0678",	x"0615",	x"0686",	
												x"302f",	x"0129",	x"0627",	x"0623",	
												x"0635",	x"0621",	x"063f",	x"062c",	
												x"062b",	x"0630",	x"061c",	x"0609",	
												x"0616",	x"0613",	x"0611",	x"0604",	
												x"0625",	x"0622",	x"065e",	x"0625",	
												x"0662",	x"0632",	x"0663",	x"063a",	
												x"0671",	x"0675",	x"0651",	x"065b",	
												x"064f",	x"0658",	x"0675",	x"064b",	
												x"0655",	x"064f",	x"0660",	x"0654",	
												x"066b",	x"0656",	x"0666",	x"064f",	
												x"0669",	x"0679",	x"068a",	x"064b",	
												x"0684",	x"0675",	x"068b",	x"0670",	
												x"065c",	x"0666",	x"066a",	x"064f",	
												x"069a",	x"0662",	x"069e",	x"066a",	
												x"0693",	x"067c",	x"069e",	x"0679",	
												x"06a2",	x"0679",	x"069e",	x"0698",	
												x"0654",	x"0685",	x"0004",	x"000a",	
												x"d441",	x"bcff",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"012a",	
												x"0644",	x"0640",	x"064b",	x"0646",	
												x"0648",	x"063f",	x"063d",	x"0625",	
												x"0639",	x"060b",	x"064e",	x"0657",	
												x"064b",	x"061b",	x"064a",	x"0630",	
												x"0681",	x"0654",	x"0686",	x"068d",	
												x"0686",	x"0666",	x"0673",	x"068d",	
												x"0684",	x"0654",	x"068b",	x"068c",	
												x"068d",	x"067b",	x"0689",	x"066b",	
												x"06b2",	x"0676",	x"06bd",	x"06bf",	
												x"06b3",	x"06c1",	x"06c9",	x"06af",	
												x"06cd",	x"06a8",	x"06b4",	x"06a4",	
												x"06aa",	x"06a9",	x"0695",	x"06a7",	
												x"06cb",	x"0694",	x"06cf",	x"06a8",	
												x"06dd",	x"06aa",	x"06ca",	x"06d6",	
												x"06cf",	x"069c",	x"06dd",	x"06bf",	
												x"06c3",	x"06be",	x"0669",	x"06b0",	
												x"502f",	x"012a",	x"0684",	x"066c",	
												x"067d",	x"068a",	x"0689",	x"0683",	
												x"068f",	x"066f",	x"0683",	x"0663",	
												x"067c",	x"0669",	x"0685",	x"0682",	
												x"067c",	x"066b",	x"06b5",	x"065f",	
												x"06c1",	x"06c1",	x"06ba",	x"06b9",	
												x"06cd",	x"06a0",	x"06c1",	x"06b7",	
												x"06cf",	x"06b6",	x"06d9",	x"06b7",	
												x"06bc",	x"06a0",	x"06d0",	x"06a0",	
												x"06d0",	x"06b3",	x"06c6",	x"06af",	
												x"06f5",	x"06b9",	x"06e2",	x"06be",	
												x"06eb",	x"06b2",	x"06e5",	x"06d5",	
												x"06c9",	x"06c4",	x"070b",	x"06b9",	
												x"070c",	x"06c8",	x"070c",	x"06eb",	
												x"070f",	x"06d3",	x"070c",	x"06e1",	
												x"071e",	x"06dc",	x"06dd",	x"06e7",	
												x"067e",	x"06c6",	x"602f",	x"012a",	
												x"068b",	x"0646",	x"06ad",	x"065a",	
												x"0690",	x"0697",	x"067b",	x"067e",	
												x"06ae",	x"065f",	x"06a1",	x"067e",	
												x"068c",	x"065f",	x"069a",	x"0667",	
												x"06d3",	x"0679",	x"06c3",	x"069f",	
												x"06df",	x"06ac",	x"06db",	x"06da",	
												x"0708",	x"06e2",	x"0702",	x"06ec",	
												x"06ef",	x"06c7",	x"06f1",	x"06e6",	
												x"06ef",	x"06e3",	x"06f5",	x"06e8",	
												x"0704",	x"06d4",	x"0720",	x"06f5",	
												x"071d",	x"06e0",	x"0731",	x"06f3",	
												x"0738",	x"06f2",	x"06fd",	x"06fc",	
												x"0711",	x"06e9",	x"0719",	x"06ed",	
												x"0727",	x"06e6",	x"0726",	x"06f1",	
												x"074e",	x"0703",	x"074e",	x"0706",	
												x"0729",	x"0709",	x"068e",	x"06f5",	
												x"702f",	x"012a",	x"06b5",	x"0660",	
												x"0703",	x"0686",	x"06a3",	x"06b3",	
												x"06c8",	x"0692",	x"06fb",	x"0686",	
												x"06fd",	x"0693",	x"06ea",	x"0697",	
												x"06af",	x"06a4",	x"0715",	x"0683",	
												x"0769",	x"06e9",	x"072f",	x"071b",	
												x"075a",	x"06f6",	x"073a",	x"06f0",	
												x"074a",	x"0713",	x"076c",	x"071b",	
												x"0722",	x"0725",	x"0760",	x"071b",	
												x"0757",	x"0727",	x"076a",	x"0727",	
												x"07a4",	x"072e",	x"0760",	x"0722",	
												x"0748",	x"074b",	x"0760",	x"072b",	
												x"0748",	x"072f",	x"0770",	x"073e",	
												x"078a",	x"074c",	x"078b",	x"0748",	
												x"07cd",	x"0771",	x"079c",	x"0794",	
												x"07b6",	x"078e",	x"0779",	x"0777",	
												x"075a",	x"0756",	x"0004",	x"000a",	
												x"1019",	x"e723",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"112b",	
												x"077a",	x"0756",	x"0792",	x"0767",	
												x"075e",	x"0772",	x"075c",	x"076f",	
												x"074b",	x"074c",	x"0741",	x"0759",	
												x"0713",	x"0725",	x"06ee",	x"06f4",	
												x"06fb",	x"06f3",	x"071f",	x"06f2",	
												x"074e",	x"0725",	x"074c",	x"074a",	
												x"0765",	x"075a",	x"0782",	x"077a",	
												x"0755",	x"0784",	x"0740",	x"076f",	
												x"074a",	x"0739",	x"075a",	x"0751",	
												x"0760",	x"0757",	x"0761",	x"0769",	
												x"0768",	x"0757",	x"0759",	x"0782",	
												x"0763",	x"075f",	x"072e",	x"0785",	
												x"074c",	x"0747",	x"074e",	x"075a",	
												x"0766",	x"0754",	x"078f",	x"0778",	
												x"075e",	x"0742",	x"0776",	x"075a",	
												x"077d",	x"0765",	x"0738",	x"0759",	
												x"102f",	x"112b",	x"072f",	x"0733",	
												x"0774",	x"073d",	x"0752",	x"075f",	
												x"074b",	x"073c",	x"0751",	x"072d",	
												x"06fc",	x"0738",	x"0703",	x"0704",	
												x"06ef",	x"06fc",	x"06d3",	x"06e2",	
												x"0707",	x"06e7",	x"0725",	x"0705",	
												x"072c",	x"0745",	x"0734",	x"0729",	
												x"075f",	x"073d",	x"0760",	x"0765",	
												x"0735",	x"0757",	x"0745",	x"0737",	
												x"0751",	x"0745",	x"074e",	x"073c",	
												x"0753",	x"074f",	x"0732",	x"075b",	
												x"0740",	x"073b",	x"074f",	x"073d",	
												x"0734",	x"0763",	x"0753",	x"0752",	
												x"074e",	x"0740",	x"0757",	x"0741",	
												x"0764",	x"075d",	x"075e",	x"0759",	
												x"076d",	x"0759",	x"076e",	x"074f",	
												x"0702",	x"075a",	x"202f",	x"112b",	
												x"0738",	x"070f",	x"072c",	x"071c",	
												x"071f",	x"0745",	x"071d",	x"0733",	
												x"06fd",	x"0719",	x"0704",	x"06f0",	
												x"06d4",	x"070e",	x"06b2",	x"06de",	
												x"06dd",	x"06de",	x"071d",	x"070b",	
												x"0711",	x"070e",	x"06fd",	x"070a",	
												x"0726",	x"0708",	x"071f",	x"073e",	
												x"0724",	x"070c",	x"06f7",	x"072a",	
												x"0737",	x"0709",	x"0757",	x"0748",	
												x"072f",	x"0730",	x"071f",	x"0742",	
												x"074c",	x"0715",	x"0755",	x"0742",	
												x"0741",	x"0739",	x"070b",	x"073d",	
												x"0738",	x"072d",	x"072d",	x"072f",	
												x"0723",	x"0730",	x"073b",	x"0737",	
												x"0756",	x"071e",	x"0750",	x"0731",	
												x"0755",	x"0747",	x"06f3",	x"0750",	
												x"302f",	x"112b",	x"0728",	x"06f9",	
												x"0715",	x"06ef",	x"072a",	x"06ec",	
												x"070c",	x"0719",	x"0706",	x"06ed",	
												x"06f6",	x"06f5",	x"070b",	x"06f1",	
												x"06de",	x"06df",	x"06e2",	x"06b8",	
												x"06e1",	x"070e",	x"0712",	x"06cc",	
												x"0721",	x"0710",	x"071b",	x"0707",	
												x"0757",	x"0740",	x"071a",	x"0762",	
												x"0720",	x"070d",	x"0729",	x"06fa",	
												x"0727",	x"0726",	x"072d",	x"071b",	
												x"0754",	x"0741",	x"074e",	x"0743",	
												x"0752",	x"0740",	x"0750",	x"073d",	
												x"071b",	x"0724",	x"074d",	x"070f",	
												x"0744",	x"0726",	x"073d",	x"0715",	
												x"0762",	x"072f",	x"0768",	x"0732",	
												x"0772",	x"073a",	x"0773",	x"0730",	
												x"070c",	x"074f",	x"0004",	x"000a",	
												x"3ae7",	x"6156",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"112c",	
												x"0714",	x"06ee",	x"0739",	x"0715",	
												x"0730",	x"070e",	x"070d",	x"0711",	
												x"073d",	x"06fe",	x"072a",	x"06fb",	
												x"0705",	x"06fc",	x"06e7",	x"06ca",	
												x"0714",	x"06d3",	x"071b",	x"06e4",	
												x"072e",	x"071b",	x"076b",	x"0712",	
												x"0763",	x"0724",	x"075e",	x"0765",	
												x"0760",	x"074d",	x"0747",	x"075b",	
												x"0779",	x"074a",	x"0777",	x"075c",	
												x"0789",	x"0770",	x"0775",	x"076b",	
												x"078c",	x"076b",	x"07a1",	x"0754",	
												x"0772",	x"0773",	x"0769",	x"0751",	
												x"0787",	x"0758",	x"0783",	x"0764",	
												x"0785",	x"076b",	x"07bb",	x"0779",	
												x"079e",	x"075b",	x"07b2",	x"0773",	
												x"07a1",	x"0787",	x"0746",	x"0782",	
												x"502f",	x"112c",	x"0757",	x"0721",	
												x"0758",	x"074e",	x"0757",	x"074c",	
												x"0756",	x"0757",	x"0744",	x"0723",	
												x"074a",	x"073e",	x"0751",	x"0730",	
												x"0723",	x"0719",	x"0759",	x"070a",	
												x"0774",	x"073f",	x"0779",	x"0752",	
												x"0792",	x"0760",	x"07a1",	x"0770",	
												x"0792",	x"077d",	x"0799",	x"0782",	
												x"079f",	x"0772",	x"0792",	x"0741",	
												x"07a4",	x"0772",	x"07ab",	x"078d",	
												x"07c4",	x"079c",	x"07d1",	x"07b9",	
												x"07ce",	x"0769",	x"07b5",	x"0779",	
												x"079a",	x"0786",	x"07bf",	x"0776",	
												x"07cf",	x"0781",	x"07cc",	x"077d",	
												x"07db",	x"077e",	x"07d4",	x"0790",	
												x"07c8",	x"0786",	x"07cf",	x"078b",	
												x"074e",	x"07aa",	x"602f",	x"112c",	
												x"0762",	x"0704",	x"0768",	x"0728",	
												x"0778",	x"0727",	x"0771",	x"071e",	
												x"077e",	x"072d",	x"0787",	x"0758",	
												x"0747",	x"0717",	x"072c",	x"0719",	
												x"0767",	x"06e3",	x"07a4",	x"06f2",	
												x"07b0",	x"0706",	x"07dd",	x"078b",	
												x"07cc",	x"077b",	x"07ce",	x"0788",	
												x"07b1",	x"07a2",	x"07bb",	x"07a7",	
												x"07c5",	x"0788",	x"080b",	x"07cb",	
												x"07d9",	x"0798",	x"07fe",	x"078b",	
												x"07f0",	x"07cd",	x"0801",	x"07c5",	
												x"07e1",	x"07ca",	x"07e6",	x"079b",	
												x"07fc",	x"07b2",	x"0811",	x"07b6",	
												x"07fb",	x"07c8",	x"0806",	x"07bc",	
												x"0829",	x"07bf",	x"0819",	x"07ba",	
												x"080b",	x"07c2",	x"077e",	x"07a9",	
												x"702f",	x"112c",	x"07a1",	x"0738",	
												x"07c1",	x"0774",	x"07b4",	x"0772",	
												x"07cf",	x"07aa",	x"07d9",	x"0761",	
												x"0763",	x"0756",	x"0788",	x"0768",	
												x"0770",	x"075f",	x"07ca",	x"0744",	
												x"07b6",	x"0764",	x"07d6",	x"076e",	
												x"0802",	x"07a3",	x"080b",	x"07cc",	
												x"0816",	x"07df",	x"081c",	x"07d1",	
												x"0804",	x"07f9",	x"0837",	x"07be",	
												x"0830",	x"07f0",	x"0845",	x"07de",	
												x"0851",	x"07f4",	x"0835",	x"0811",	
												x"0847",	x"0807",	x"0860",	x"0817",	
												x"07fd",	x"0819",	x"0864",	x"080d",	
												x"0874",	x"0842",	x"084f",	x"083e",	
												x"084d",	x"0845",	x"088e",	x"0820",	
												x"086b",	x"084b",	x"0870",	x"083c",	
												x"06f5",	x"084f",	x"0004",	x"000a",	
												x"7599",	x"85fc",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"212d",	
												x"0707",	x"0705",	x"06ec",	x"0707",	
												x"06ee",	x"06f5",	x"06f9",	x"06db",	
												x"06da",	x"06e7",	x"06b9",	x"06bc",	
												x"06c9",	x"06d0",	x"068f",	x"06bc",	
												x"06b0",	x"06a6",	x"06cb",	x"06ba",	
												x"06cc",	x"06d8",	x"0700",	x"0703",	
												x"06f9",	x"06f2",	x"071c",	x"06e0",	
												x"06f3",	x"070c",	x"06c4",	x"06f7",	
												x"06f7",	x"06eb",	x"06f9",	x"0711",	
												x"0709",	x"06ee",	x"06ff",	x"06f0",	
												x"0705",	x"06e6",	x"06fd",	x"0702",	
												x"0704",	x"06fc",	x"06b6",	x"06fe",	
												x"0706",	x"06c4",	x"071b",	x"0709",	
												x"0725",	x"0719",	x"0711",	x"06fd",	
												x"0708",	x"0713",	x"0731",	x"0707",	
												x"0730",	x"0720",	x"06aa",	x"0715",	
												x"102f",	x"212d",	x"06c7",	x"06ba",	
												x"06ca",	x"06e1",	x"06fc",	x"06de",	
												x"06fc",	x"06e1",	x"06d2",	x"06cb",	
												x"06a9",	x"06ab",	x"0687",	x"068a",	
												x"065f",	x"067f",	x"06bb",	x"066b",	
												x"06da",	x"06ad",	x"06e5",	x"06b1",	
												x"06f5",	x"06d2",	x"06f9",	x"06fa",	
												x"0703",	x"06fe",	x"06d1",	x"0712",	
												x"06cd",	x"06f8",	x"06d8",	x"06c1",	
												x"06eb",	x"06e3",	x"06fb",	x"06e6",	
												x"06f7",	x"0705",	x"06f3",	x"0710",	
												x"0711",	x"0708",	x"0716",	x"0708",	
												x"06c9",	x"06f3",	x"06f0",	x"06eb",	
												x"06f2",	x"06fe",	x"0701",	x"06e3",	
												x"06ef",	x"0702",	x"0704",	x"06f6",	
												x"0714",	x"070e",	x"0709",	x"0701",	
												x"06be",	x"06ec",	x"202f",	x"212d",	
												x"06be",	x"06c5",	x"0694",	x"06cb",	
												x"06dd",	x"06a1",	x"06e1",	x"06e1",	
												x"06b4",	x"06d0",	x"0684",	x"06aa",	
												x"0680",	x"066d",	x"0635",	x"067d",	
												x"06b2",	x"066f",	x"06b2",	x"06cf",	
												x"06cd",	x"06cc",	x"06cc",	x"06e5",	
												x"06de",	x"06c3",	x"0701",	x"06db",	
												x"06d6",	x"06db",	x"06be",	x"06d8",	
												x"06cc",	x"06c5",	x"06d8",	x"06ce",	
												x"06d6",	x"06c3",	x"06e1",	x"06d4",	
												x"06c6",	x"06db",	x"06f7",	x"06dc",	
												x"06d5",	x"06de",	x"06d3",	x"06c9",	
												x"06e2",	x"06d8",	x"06df",	x"06d9",	
												x"06d5",	x"06c8",	x"06e4",	x"06eb",	
												x"06f7",	x"06c8",	x"0713",	x"06ea",	
												x"0702",	x"06f3",	x"06a6",	x"06ef",	
												x"302f",	x"212d",	x"06a4",	x"069c",	
												x"06c5",	x"069e",	x"06af",	x"069e",	
												x"06d7",	x"0698",	x"06bd",	x"0696",	
												x"0690",	x"0689",	x"0689",	x"0692",	
												x"068c",	x"066e",	x"06aa",	x"066b",	
												x"06ba",	x"0694",	x"06cb",	x"06bd",	
												x"06d0",	x"06aa",	x"06d2",	x"06ab",	
												x"06ed",	x"06d1",	x"06d7",	x"06c9",	
												x"06ab",	x"06bb",	x"06da",	x"069c",	
												x"06e9",	x"06c9",	x"06f3",	x"06cf",	
												x"06e6",	x"06cf",	x"06ee",	x"06d3",	
												x"06fa",	x"0706",	x"0702",	x"06e4",	
												x"06bc",	x"06d8",	x"0718",	x"06da",	
												x"06de",	x"06ed",	x"06e4",	x"06d4",	
												x"06ee",	x"06cb",	x"0724",	x"06ce",	
												x"0722",	x"06fc",	x"0726",	x"06fd",	
												x"069f",	x"06f6",	x"0004",	x"000a",	
												x"0dc9",	x"7369",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"212e",	
												x"06ce",	x"0697",	x"06e5",	x"06b6",	
												x"06e0",	x"06c6",	x"06e3",	x"06d9",	
												x"06ca",	x"06cc",	x"0699",	x"06a6",	
												x"06a3",	x"069e",	x"0685",	x"0691",	
												x"06c6",	x"0695",	x"06e7",	x"06c8",	
												x"0713",	x"06dc",	x"0723",	x"071f",	
												x"0706",	x"06e7",	x"06fb",	x"0700",	
												x"06ff",	x"070a",	x"06f5",	x"070f",	
												x"0709",	x"06fa",	x"071d",	x"071f",	
												x"0733",	x"070b",	x"0721",	x"071c",	
												x"0737",	x"0728",	x"072d",	x"0715",	
												x"073e",	x"0719",	x"070d",	x"070e",	
												x"0742",	x"0708",	x"072f",	x"073d",	
												x"073f",	x"070e",	x"075d",	x"0727",	
												x"076c",	x"0726",	x"0774",	x"0747",	
												x"076b",	x"072f",	x"06dc",	x"071c",	
												x"502f",	x"212e",	x"0713",	x"06db",	
												x"070d",	x"06fc",	x"0718",	x"06e5",	
												x"071a",	x"0722",	x"06eb",	x"06c5",	
												x"06e7",	x"06d2",	x"06ee",	x"06bc",	
												x"06c3",	x"06bd",	x"071f",	x"06af",	
												x"0741",	x"0714",	x"0715",	x"0707",	
												x"0753",	x"072b",	x"074e",	x"0725",	
												x"0757",	x"074a",	x"0761",	x"0727",	
												x"071e",	x"072e",	x"0752",	x"070e",	
												x"074d",	x"074b",	x"0751",	x"071d",	
												x"076e",	x"0744",	x"076c",	x"074a",	
												x"0776",	x"073f",	x"0762",	x"0736",	
												x"073b",	x"0735",	x"076c",	x"0731",	
												x"0751",	x"0743",	x"076a",	x"071d",	
												x"077d",	x"0734",	x"0792",	x"073d",	
												x"0794",	x"0747",	x"0799",	x"0741",	
												x"070b",	x"0747",	x"602f",	x"212e",	
												x"06fe",	x"06cc",	x"070d",	x"06ea",	
												x"06fe",	x"06ac",	x"0701",	x"06e7",	
												x"0716",	x"06ea",	x"072a",	x"06c8",	
												x"0716",	x"06a0",	x"0713",	x"06d0",	
												x"0755",	x"06cd",	x"074a",	x"070a",	
												x"0743",	x"0715",	x"078a",	x"072f",	
												x"0794",	x"0744",	x"0776",	x"0753",	
												x"0768",	x"072f",	x"076c",	x"0741",	
												x"0783",	x"0744",	x"078f",	x"076a",	
												x"077c",	x"072f",	x"07a1",	x"075a",	
												x"0799",	x"0767",	x"07a0",	x"0766",	
												x"0784",	x"0755",	x"078c",	x"0742",	
												x"079f",	x"075e",	x"078a",	x"074b",	
												x"07ad",	x"0757",	x"07b4",	x"076d",	
												x"07cf",	x"076a",	x"07d0",	x"0773",	
												x"07ca",	x"077d",	x"070f",	x"0792",	
												x"702f",	x"212e",	x"072a",	x"06e8",	
												x"073f",	x"070e",	x"075f",	x"0715",	
												x"0748",	x"0721",	x"0725",	x"070e",	
												x"073c",	x"0730",	x"073b",	x"06d4",	
												x"071a",	x"06e0",	x"07aa",	x"06ee",	
												x"0786",	x"06fb",	x"0791",	x"0739",	
												x"07a7",	x"0772",	x"07a5",	x"077b",	
												x"07c2",	x"0774",	x"07c1",	x"07b5",	
												x"07ad",	x"076e",	x"07f1",	x"07a2",	
												x"07de",	x"078f",	x"07ee",	x"078e",	
												x"07ed",	x"07a0",	x"0806",	x"07c5",	
												x"07ed",	x"07d3",	x"080e",	x"07b6",	
												x"07cf",	x"07b7",	x"07f1",	x"079e",	
												x"07e1",	x"07ca",	x"07f0",	x"07a3",	
												x"07f9",	x"07d1",	x"082c",	x"07cb",	
												x"0843",	x"07d7",	x"0813",	x"0809",	
												x"0711",	x"07e2",	x"0004",	x"000a",	
												x"4bdc",	x"9e9b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"312f",	
												x"073a",	x"072f",	x"073f",	x"0748",	
												x"0752",	x"0738",	x"074a",	x"074a",	
												x"0723",	x"072e",	x"0735",	x"0712",	
												x"0730",	x"071d",	x"06dd",	x"06e5",	
												x"06f6",	x"06d2",	x"0717",	x"070f",	
												x"071b",	x"071f",	x"0737",	x"072c",	
												x"0723",	x"075b",	x"073e",	x"0757",	
												x"0758",	x"0747",	x"0725",	x"075d",	
												x"073e",	x"072a",	x"0764",	x"0769",	
												x"0733",	x"074b",	x"0760",	x"0752",	
												x"072d",	x"0739",	x"073b",	x"0739",	
												x"073a",	x"0755",	x"0734",	x"0729",	
												x"0756",	x"0759",	x"073c",	x"075c",	
												x"0744",	x"072d",	x"0746",	x"0746",	
												x"0756",	x"0733",	x"0754",	x"0752",	
												x"0743",	x"0729",	x"0711",	x"073d",	
												x"102f",	x"312f",	x"0709",	x"06f7",	
												x"073a",	x"0742",	x"0711",	x"0735",	
												x"071d",	x"072d",	x"06f4",	x"06f8",	
												x"0701",	x"06f6",	x"06ee",	x"06ef",	
												x"06ad",	x"06f0",	x"0701",	x"069c",	
												x"0705",	x"06e9",	x"0702",	x"070d",	
												x"0712",	x"0713",	x"072d",	x"072f",	
												x"073e",	x"0751",	x"0727",	x"0750",	
												x"06dd",	x"0738",	x"0716",	x"0740",	
												x"0739",	x"0751",	x"0722",	x"072f",	
												x"074c",	x"072c",	x"072e",	x"073b",	
												x"0732",	x"073d",	x"0746",	x"0739",	
												x"071e",	x"0736",	x"073e",	x"074a",	
												x"0734",	x"072d",	x"0726",	x"072b",	
												x"0736",	x"0732",	x"072a",	x"071b",	
												x"073e",	x"073a",	x"076b",	x"0752",	
												x"06d2",	x"074d",	x"202f",	x"312f",	
												x"06f0",	x"06e6",	x"06f7",	x"071f",	
												x"0713",	x"0714",	x"06f8",	x"0711",	
												x"06f4",	x"06ef",	x"06d6",	x"06f7",	
												x"06d1",	x"06ed",	x"06b0",	x"06f6",	
												x"06c4",	x"0697",	x"06ee",	x"06e6",	
												x"0704",	x"0721",	x"06fe",	x"06fb",	
												x"0709",	x"06fa",	x"06ea",	x"072c",	
												x"073e",	x"06fd",	x"06ed",	x"0728",	
												x"0714",	x"0704",	x"0718",	x"0714",	
												x"06fa",	x"072c",	x"071e",	x"06fd",	
												x"0728",	x"071e",	x"0727",	x"0720",	
												x"0719",	x"0714",	x"072e",	x"071f",	
												x"074e",	x"071d",	x"072b",	x"072d",	
												x"0720",	x"0737",	x"072c",	x"0714",	
												x"0725",	x"0722",	x"0757",	x"071c",	
												x"0748",	x"0716",	x"06c6",	x"0712",	
												x"302f",	x"312f",	x"06e3",	x"06cb",	
												x"06f1",	x"06d6",	x"06f8",	x"06d9",	
												x"06ea",	x"06e4",	x"06f6",	x"06cf",	
												x"06f4",	x"06ce",	x"06a7",	x"06b7",	
												x"0695",	x"06b8",	x"06e8",	x"068b",	
												x"06e8",	x"06df",	x"06fc",	x"06d8",	
												x"0702",	x"06d8",	x"0712",	x"06e5",	
												x"0703",	x"0715",	x"0701",	x"06f6",	
												x"06d5",	x"0700",	x"070d",	x"06e0",	
												x"0715",	x"0710",	x"0724",	x"0711",	
												x"071d",	x"071e",	x"073c",	x"072a",	
												x"0739",	x"0735",	x"0711",	x"071b",	
												x"072c",	x"06fe",	x"073c",	x"0724",	
												x"0721",	x"072b",	x"072f",	x"06ee",	
												x"0720",	x"0716",	x"0741",	x"0700",	
												x"0757",	x"071d",	x"074e",	x"0726",	
												x"06e2",	x"071e",	x"0004",	x"000a",	
												x"2c48",	x"d48e",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"3130",	
												x"0703",	x"06e8",	x"070a",	x"0700",	
												x"070d",	x"06bb",	x"0719",	x"0708",	
												x"06f6",	x"06de",	x"06f8",	x"06ea",	
												x"06f8",	x"06ec",	x"06d0",	x"0702",	
												x"06fd",	x"06a9",	x"072f",	x"06da",	
												x"0721",	x"06e4",	x"0737",	x"0718",	
												x"0746",	x"070e",	x"0740",	x"073c",	
												x"0743",	x"0738",	x"0749",	x"0727",	
												x"075d",	x"0702",	x"077e",	x"0752",	
												x"0753",	x"075b",	x"076a",	x"0754",	
												x"076a",	x"0741",	x"075a",	x"074d",	
												x"0772",	x"0758",	x"075d",	x"0752",	
												x"0769",	x"0746",	x"0756",	x"0745",	
												x"076d",	x"074f",	x"0770",	x"0763",	
												x"0798",	x"074a",	x"0794",	x"076b",	
												x"0792",	x"0773",	x"0713",	x"0764",	
												x"502f",	x"3130",	x"071f",	x"06ef",	
												x"0750",	x"0738",	x"074b",	x"0738",	
												x"0737",	x"073f",	x"0757",	x"0715",	
												x"0735",	x"0715",	x"0720",	x"071d",	
												x"070b",	x"06f5",	x"0767",	x"06fc",	
												x"0768",	x"0717",	x"0789",	x"072a",	
												x"0783",	x"075e",	x"0789",	x"073f",	
												x"07ad",	x"074b",	x"0792",	x"0745",	
												x"075e",	x"0732",	x"07a5",	x"074a",	
												x"0795",	x"077f",	x"078c",	x"0747",	
												x"079b",	x"0789",	x"078f",	x"0765",	
												x"0793",	x"0769",	x"079d",	x"0761",	
												x"079c",	x"0750",	x"07bc",	x"077c",	
												x"07be",	x"076e",	x"07c3",	x"0757",	
												x"07cd",	x"0780",	x"07a8",	x"0772",	
												x"07f3",	x"078f",	x"07c0",	x"0790",	
												x"0727",	x"078f",	x"602f",	x"3130",	
												x"075e",	x"06fa",	x"0756",	x"070f",	
												x"0772",	x"0725",	x"0750",	x"0755",	
												x"0744",	x"071f",	x"0740",	x"072c",	
												x"0731",	x"070b",	x"0736",	x"06eb",	
												x"076f",	x"0700",	x"077e",	x"06fc",	
												x"079c",	x"0744",	x"07ba",	x"0748",	
												x"07ae",	x"0786",	x"078b",	x"0780",	
												x"07a5",	x"076e",	x"077d",	x"077a",	
												x"07b9",	x"076b",	x"07a5",	x"078f",	
												x"07b1",	x"0792",	x"07f9",	x"07a6",	
												x"07ba",	x"0780",	x"07e4",	x"0797",	
												x"07ce",	x"079f",	x"07bd",	x"07af",	
												x"07d1",	x"0793",	x"07e0",	x"07ba",	
												x"07dd",	x"078e",	x"07fd",	x"07aa",	
												x"07fd",	x"0796",	x"07ed",	x"07a1",	
												x"082b",	x"07a6",	x"0743",	x"079f",	
												x"702f",	x"3130",	x"0799",	x"0723",	
												x"079e",	x"076f",	x"0780",	x"0787",	
												x"07c2",	x"076d",	x"0774",	x"073c",	
												x"0771",	x"074e",	x"077f",	x"074a",	
												x"0771",	x"0755",	x"07c5",	x"073f",	
												x"07a7",	x"074a",	x"07ef",	x"0765",	
												x"0826",	x"079a",	x"07f6",	x"07ba",	
												x"07ee",	x"07a8",	x"07fb",	x"07a3",	
												x"0801",	x"07d4",	x"080c",	x"07da",	
												x"080d",	x"07db",	x"0829",	x"07d6",	
												x"084e",	x"07f5",	x"0828",	x"07e1",	
												x"084c",	x"07ff",	x"082e",	x"0811",	
												x"082c",	x"081a",	x"083b",	x"07f0",	
												x"0850",	x"07fa",	x"0842",	x"07fd",	
												x"0859",	x"0811",	x"0862",	x"0815",	
												x"0874",	x"0833",	x"088c",	x"083a",	
												x"065d",	x"0823",	x"0004",	x"000a",	
												x"69a5",	x"fab6",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"0131",	
												x"066a",	x"068f",	x"065a",	x"0656",	
												x"065a",	x"0663",	x"0645",	x"0662",	
												x"0659",	x"0638",	x"068b",	x"0642",	
												x"069f",	x"0695",	x"0655",	x"06d2",	
												x"068c",	x"0664",	x"06bb",	x"06bd",	
												x"06b0",	x"06b0",	x"0690",	x"0696",	
												x"0692",	x"0694",	x"0682",	x"068c",	
												x"0694",	x"068a",	x"062a",	x"068d",	
												x"0666",	x"065b",	x"0699",	x"0696",	
												x"068a",	x"0691",	x"0695",	x"0693",	
												x"06a0",	x"069b",	x"069a",	x"068e",	
												x"069e",	x"06b5",	x"0661",	x"0698",	
												x"0687",	x"0667",	x"06a9",	x"06af",	
												x"06a5",	x"06ab",	x"069f",	x"06b2",	
												x"06a7",	x"069c",	x"06d1",	x"0697",	
												x"0691",	x"06a0",	x"064a",	x"0681",	
												x"1030",	x"0131",	x"0637",	x"065a",	
												x"0631",	x"063a",	x"0634",	x"0631",	
												x"061c",	x"065e",	x"0656",	x"0621",	
												x"067b",	x"063e",	x"0679",	x"0660",	
												x"064b",	x"0672",	x"0647",	x"066f",	
												x"0685",	x"067d",	x"0685",	x"068c",	
												x"0655",	x"0686",	x"0680",	x"068d",	
												x"0695",	x"069f",	x"068f",	x"06a3",	
												x"0615",	x"069e",	x"0673",	x"0668",	
												x"066e",	x"068e",	x"065b",	x"0672",	
												x"0681",	x"0689",	x"068f",	x"0679",	
												x"067c",	x"068a",	x"0674",	x"0675",	
												x"0644",	x"0691",	x"0678",	x"0687",	
												x"067c",	x"0691",	x"068b",	x"0690",	
												x"068c",	x"0687",	x"0690",	x"068f",	
												x"0697",	x"06b0",	x"067e",	x"0697",	
												x"0637",	x"0679",	x"2030",	x"0131",	
												x"0647",	x"064c",	x"0657",	x"063c",	
												x"0607",	x"0645",	x"0618",	x"061e",	
												x"0629",	x"0644",	x"0665",	x"0673",	
												x"064f",	x"067f",	x"063a",	x"066d",	
												x"063e",	x"064f",	x"063d",	x"0656",	
												x"064d",	x"0660",	x"065e",	x"0651",	
												x"0664",	x"067e",	x"0669",	x"0674",	
												x"0659",	x"066a",	x"063f",	x"0675",	
												x"065d",	x"0665",	x"064e",	x"065e",	
												x"0643",	x"064c",	x"0647",	x"066e",	
												x"064d",	x"0663",	x"0681",	x"064b",	
												x"0677",	x"0687",	x"0639",	x"0656",	
												x"0670",	x"0653",	x"0672",	x"066b",	
												x"0673",	x"067a",	x"0681",	x"067d",	
												x"064b",	x"066c",	x"0685",	x"0665",	
												x"065d",	x"0663",	x"062d",	x"065e",	
												x"3030",	x"0131",	x"063e",	x"0634",	
												x"061b",	x"0615",	x"061c",	x"0607",	
												x"0618",	x"0621",	x"0632",	x"0609",	
												x"0654",	x"0638",	x"064f",	x"0650",	
												x"061e",	x"0645",	x"0636",	x"063b",	
												x"065c",	x"0644",	x"065c",	x"064d",	
												x"0659",	x"0666",	x"0657",	x"0659",	
												x"067c",	x"0662",	x"0660",	x"066d",	
												x"0628",	x"0655",	x"063d",	x"0632",	
												x"0649",	x"064b",	x"063e",	x"0653",	
												x"065e",	x"0655",	x"0674",	x"065b",	
												x"0691",	x"0676",	x"066b",	x"0682",	
												x"0622",	x"065b",	x"066e",	x"0642",	
												x"067f",	x"066f",	x"067a",	x"0660",	
												x"0691",	x"0670",	x"0699",	x"066b",	
												x"0695",	x"0676",	x"0680",	x"0665",	
												x"0628",	x"0682",	x"0004",	x"000a",	
												x"d247",	x"bf7a",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"0132",	
												x"063a",	x"064d",	x"0629",	x"0632",	
												x"0620",	x"0600",	x"0634",	x"0622",	
												x"062f",	x"060d",	x"0659",	x"064f",	
												x"066f",	x"0665",	x"064d",	x"0640",	
												x"0671",	x"063d",	x"066b",	x"065e",	
												x"0681",	x"065b",	x"0678",	x"069b",	
												x"067b",	x"0662",	x"0689",	x"067c",	
												x"068d",	x"0691",	x"0649",	x"0689",	
												x"069c",	x"0650",	x"067e",	x"0668",	
												x"0686",	x"0697",	x"0693",	x"067f",	
												x"06a0",	x"06a0",	x"069c",	x"069b",	
												x"0687",	x"069e",	x"0676",	x"0696",	
												x"0697",	x"0686",	x"06b7",	x"0698",	
												x"06b7",	x"06a1",	x"06bc",	x"06bd",	
												x"06be",	x"069d",	x"06ba",	x"06b4",	
												x"06b3",	x"06a7",	x"067a",	x"06ba",	
												x"5030",	x"0132",	x"0670",	x"066e",	
												x"0667",	x"065d",	x"0663",	x"064c",	
												x"068a",	x"0678",	x"068a",	x"0684",	
												x"0685",	x"0683",	x"068f",	x"068a",	
												x"0687",	x"0696",	x"0698",	x"0684",	
												x"06be",	x"0692",	x"06a8",	x"0691",	
												x"06be",	x"06a2",	x"06b8",	x"06b8",	
												x"06b7",	x"06b7",	x"06b7",	x"06b5",	
												x"06b2",	x"069f",	x"06a7",	x"068c",	
												x"06a9",	x"06aa",	x"06b1",	x"069e",	
												x"06c0",	x"06b8",	x"06d4",	x"06b9",	
												x"06c0",	x"06b0",	x"06b2",	x"06b1",	
												x"06a6",	x"069e",	x"06e8",	x"06a5",	
												x"06c9",	x"06bb",	x"06f0",	x"06cb",	
												x"0704",	x"06cd",	x"06e8",	x"06c5",	
												x"06e9",	x"06ba",	x"06cd",	x"06cf",	
												x"0693",	x"06c0",	x"6030",	x"0132",	
												x"06a0",	x"0697",	x"0690",	x"0674",	
												x"0692",	x"067b",	x"06a0",	x"0684",	
												x"06af",	x"0675",	x"0697",	x"0694",	
												x"069f",	x"0694",	x"069f",	x"06a1",	
												x"0699",	x"067c",	x"06ec",	x"0681",	
												x"06be",	x"06c2",	x"06e6",	x"06c9",	
												x"06f8",	x"06e6",	x"06db",	x"06e0",	
												x"06d0",	x"06e7",	x"06cc",	x"06cb",	
												x"06e1",	x"06b2",	x"06d8",	x"06cf",	
												x"06ef",	x"06d4",	x"0709",	x"06ec",	
												x"0703",	x"06e9",	x"070c",	x"06ea",	
												x"06fc",	x"06fe",	x"06d0",	x"06c9",	
												x"0714",	x"06d0",	x"070c",	x"0704",	
												x"070c",	x"0700",	x"0718",	x"06fe",	
												x"0716",	x"06f6",	x"073a",	x"06f0",	
												x"072f",	x"06f8",	x"06d5",	x"070a",	
												x"7030",	x"0132",	x"070b",	x"06c1",	
												x"06c6",	x"0685",	x"069f",	x"068e",	
												x"06d9",	x"06a5",	x"06e2",	x"06bb",	
												x"0708",	x"06e2",	x"06ee",	x"06f9",	
												x"06d7",	x"06bd",	x"0723",	x"06d3",	
												x"072b",	x"0719",	x"0718",	x"0721",	
												x"0746",	x"0715",	x"0765",	x"072c",	
												x"075b",	x"0748",	x"0739",	x"073b",	
												x"0704",	x"073a",	x"0743",	x"0708",	
												x"0733",	x"073e",	x"074a",	x"0722",	
												x"0778",	x"0742",	x"0787",	x"076f",	
												x"077b",	x"077b",	x"0746",	x"076e",	
												x"0744",	x"075f",	x"076f",	x"0760",	
												x"079c",	x"0770",	x"0780",	x"0771",	
												x"07b5",	x"0793",	x"07a1",	x"077a",	
												x"07b4",	x"077b",	x"0781",	x"0788",	
												x"0720",	x"0779",	x"0004",	x"000a",	
												x"0855",	x"e939",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"1133",	
												x"0709",	x"0745",	x"0716",	x"06ee",	
												x"0705",	x"0722",	x"0707",	x"072a",	
												x"070e",	x"06ff",	x"071a",	x"0713",	
												x"0720",	x"071f",	x"070f",	x"073d",	
												x"0764",	x"072f",	x"075f",	x"076b",	
												x"0760",	x"0770",	x"074e",	x"0771",	
												x"072e",	x"0773",	x"073f",	x"0753",	
												x"0739",	x"074b",	x"0710",	x"0776",	
												x"0733",	x"0747",	x"074c",	x"0761",	
												x"073b",	x"0751",	x"0760",	x"075d",	
												x"0746",	x"0750",	x"075d",	x"0735",	
												x"073a",	x"0754",	x"06fa",	x"0734",	
												x"075d",	x"06fc",	x"0747",	x"0752",	
												x"0752",	x"0748",	x"0769",	x"074c",	
												x"073c",	x"0744",	x"0777",	x"0761",	
												x"0749",	x"074f",	x"0718",	x"073c",	
												x"1030",	x"1133",	x"06ff",	x"06f7",	
												x"0704",	x"0720",	x"06e4",	x"0709",	
												x"06fc",	x"070b",	x"0702",	x"06e7",	
												x"0703",	x"06f7",	x"0720",	x"0710",	
												x"0707",	x"072b",	x"073c",	x"073a",	
												x"0737",	x"0737",	x"0736",	x"072e",	
												x"0735",	x"0747",	x"0737",	x"072e",	
												x"0739",	x"0734",	x"0758",	x"0753",	
												x"070d",	x"076f",	x"0720",	x"0738",	
												x"0743",	x"074c",	x"074d",	x"0745",	
												x"071b",	x"075e",	x"0732",	x"0740",	
												x"0732",	x"072d",	x"0741",	x"0725",	
												x"071e",	x"0736",	x"074d",	x"0740",	
												x"075a",	x"073f",	x"0761",	x"074e",	
												x"0755",	x"0753",	x"074f",	x"073e",	
												x"074a",	x"0754",	x"076a",	x"0730",	
												x"06e1",	x"0746",	x"2030",	x"1133",	
												x"06dd",	x"0706",	x"06e2",	x"06f6",	
												x"06f0",	x"0706",	x"06fc",	x"070d",	
												x"06fe",	x"0714",	x"071b",	x"0711",	
												x"0730",	x"0730",	x"0713",	x"073d",	
												x"0719",	x"072c",	x"0731",	x"0753",	
												x"0730",	x"072f",	x"0705",	x"071a",	
												x"0712",	x"0715",	x"0728",	x"0724",	
												x"072c",	x"0732",	x"0703",	x"0745",	
												x"071c",	x"06fe",	x"0728",	x"0726",	
												x"071e",	x"0719",	x"0716",	x"0715",	
												x"0725",	x"0711",	x"073c",	x"0736",	
												x"071e",	x"071c",	x"0705",	x"0718",	
												x"0729",	x"0717",	x"072a",	x"0755",	
												x"0741",	x"0731",	x"0751",	x"074c",	
												x"074f",	x"0737",	x"0742",	x"073c",	
												x"073d",	x"0716",	x"06e8",	x"0733",	
												x"3030",	x"1133",	x"06cf",	x"06d8",	
												x"06df",	x"06d6",	x"06dd",	x"06d8",	
												x"06f6",	x"06dc",	x"06e4",	x"06e4",	
												x"06d6",	x"06e7",	x"06fc",	x"06e4",	
												x"06cc",	x"06e1",	x"0709",	x"06ea",	
												x"072a",	x"0705",	x"072a",	x"0719",	
												x"06f2",	x"071f",	x"0712",	x"06f9",	
												x"0733",	x"0713",	x"0714",	x"072b",	
												x"0713",	x"0719",	x"0738",	x"0716",	
												x"0726",	x"0722",	x"0717",	x"071f",	
												x"0712",	x"0722",	x"0712",	x"070d",	
												x"0718",	x"0708",	x"0740",	x"071a",	
												x"071c",	x"072f",	x"074e",	x"071b",	
												x"074a",	x"075b",	x"0745",	x"073c",	
												x"0745",	x"0735",	x"074b",	x"0724",	
												x"074d",	x"0728",	x"0744",	x"0722",	
												x"06ee",	x"0727",	x"0004",	x"000a",	
												x"3277",	x"5dcb",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"1134",	
												x"06f0",	x"06fb",	x"06f8",	x"06e6",	
												x"070a",	x"06d2",	x"0709",	x"070a",	
												x"0725",	x"0700",	x"072b",	x"071c",	
												x"0723",	x"0723",	x"0702",	x"0735",	
												x"071e",	x"0704",	x"0744",	x"0718",	
												x"074b",	x"0733",	x"0755",	x"0739",	
												x"0742",	x"0741",	x"0744",	x"073f",	
												x"0743",	x"0752",	x"0732",	x"0737",	
												x"077b",	x"0740",	x"074c",	x"0749",	
												x"076b",	x"0741",	x"0749",	x"075f",	
												x"0759",	x"0744",	x"0759",	x"0752",	
												x"076f",	x"0756",	x"075e",	x"0762",	
												x"0774",	x"075b",	x"0774",	x"0768",	
												x"0779",	x"077e",	x"0788",	x"077e",	
												x"078d",	x"0779",	x"079d",	x"077b",	
												x"0783",	x"0770",	x"0730",	x"076a",	
												x"5030",	x"1134",	x"072b",	x"0738",	
												x"0728",	x"0733",	x"073e",	x"0723",	
												x"0752",	x"0725",	x"0739",	x"074c",	
												x"0776",	x"075f",	x"0751",	x"0753",	
												x"0748",	x"074d",	x"0783",	x"0748",	
												x"076f",	x"0778",	x"0765",	x"0756",	
												x"0782",	x"0774",	x"0785",	x"0781",	
												x"077a",	x"0773",	x"0762",	x"076b",	
												x"0766",	x"0754",	x"078c",	x"0756",	
												x"078b",	x"0783",	x"078a",	x"0780",	
												x"078f",	x"0779",	x"07b8",	x"076e",	
												x"07b0",	x"0779",	x"07a4",	x"0781",	
												x"079e",	x"0777",	x"079a",	x"075f",	
												x"07b1",	x"0780",	x"07af",	x"0781",	
												x"07b7",	x"0777",	x"07a3",	x"0789",	
												x"07c5",	x"077c",	x"07c4",	x"078e",	
												x"072c",	x"0797",	x"6030",	x"1134",	
												x"0749",	x"06f4",	x"074d",	x"0728",	
												x"075e",	x"073d",	x"0760",	x"0743",	
												x"0748",	x"0748",	x"0769",	x"0736",	
												x"075f",	x"077e",	x"0765",	x"0751",	
												x"0794",	x"075b",	x"07a3",	x"0789",	
												x"079e",	x"078d",	x"07a7",	x"07a6",	
												x"07b0",	x"07a8",	x"07b1",	x"079a",	
												x"07b1",	x"0775",	x"07ac",	x"079c",	
												x"07a7",	x"07a1",	x"07ba",	x"07c7",	
												x"07ae",	x"07ab",	x"07b0",	x"07bd",	
												x"07b1",	x"07a0",	x"07c5",	x"07a9",	
												x"07c3",	x"07ae",	x"07bb",	x"07b0",	
												x"07e3",	x"0787",	x"07f8",	x"07c3",	
												x"07ff",	x"07cd",	x"0800",	x"07c8",	
												x"080f",	x"07bf",	x"07ea",	x"07cf",	
												x"07d8",	x"07ca",	x"07ac",	x"07ab",	
												x"7030",	x"1134",	x"07c5",	x"078f",	
												x"07af",	x"0795",	x"07c8",	x"078a",	
												x"07dc",	x"0774",	x"07ac",	x"0785",	
												x"07d6",	x"0793",	x"07d8",	x"07bc",	
												x"07ee",	x"07d5",	x"07f4",	x"0789",	
												x"0820",	x"07ce",	x"081f",	x"07f6",	
												x"0805",	x"0807",	x"0805",	x"07f8",	
												x"0829",	x"0816",	x"081f",	x"0807",	
												x"080a",	x"0803",	x"081c",	x"07f6",	
												x"0825",	x"0821",	x"0840",	x"080d",	
												x"084a",	x"081d",	x"0845",	x"0817",	
												x"0853",	x"0830",	x"0835",	x"0832",	
												x"0835",	x"0838",	x"084b",	x"0843",	
												x"0850",	x"0848",	x"0850",	x"0857",	
												x"0862",	x"084b",	x"0879",	x"084d",	
												x"0843",	x"0843",	x"0868",	x"083b",	
												x"06da",	x"084b",	x"0004",	x"000a",	
												x"6f8b",	x"8e8b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"2135",	
												x"06a7",	x"06e4",	x"069e",	x"06a1",	
												x"06cc",	x"0699",	x"06bf",	x"06c0",	
												x"06ba",	x"06c3",	x"06ba",	x"06e6",	
												x"06ba",	x"06e0",	x"06c4",	x"06e8",	
												x"06f0",	x"06c4",	x"0701",	x"06eb",	
												x"06ec",	x"06ed",	x"06ee",	x"0709",	
												x"0700",	x"06f5",	x"0710",	x"06d3",	
												x"06f0",	x"0711",	x"06a0",	x"0702",	
												x"06dc",	x"06d5",	x"06cc",	x"0703",	
												x"072c",	x"0700",	x"06e1",	x"0702",	
												x"06fb",	x"06f2",	x"06ff",	x"0712",	
												x"06eb",	x"0702",	x"06ac",	x"06e8",	
												x"0706",	x"06e0",	x"0725",	x"070e",	
												x"0721",	x"06ff",	x"0720",	x"0718",	
												x"06f5",	x"06f8",	x"06ff",	x"06e0",	
												x"06e2",	x"06e8",	x"0677",	x"06ed",	
												x"1030",	x"2135",	x"06b8",	x"0692",	
												x"06a8",	x"06b1",	x"067f",	x"06a4",	
												x"06b1",	x"069a",	x"06c5",	x"06ab",	
												x"06dd",	x"06ca",	x"06d8",	x"06e9",	
												x"06b4",	x"06c5",	x"06f0",	x"06c3",	
												x"0706",	x"06fd",	x"070d",	x"06f6",	
												x"06e6",	x"06f7",	x"06e1",	x"06f4",	
												x"06d6",	x"06d8",	x"06c3",	x"06f8",	
												x"06a9",	x"06f3",	x"06d7",	x"06d2",	
												x"06ce",	x"06dd",	x"06e3",	x"06ee",	
												x"06e9",	x"06fb",	x"06ed",	x"06eb",	
												x"06ed",	x"06ff",	x"06e1",	x"06f1",	
												x"06a8",	x"06ec",	x"06f0",	x"06d7",	
												x"06f0",	x"06ef",	x"06f6",	x"06f1",	
												x"06ef",	x"06f9",	x"0728",	x"06ef",	
												x"06f9",	x"0707",	x"0706",	x"06fb",	
												x"0686",	x"06f2",	x"2030",	x"2135",	
												x"0685",	x"0693",	x"06a4",	x"069a",	
												x"06a2",	x"0692",	x"069b",	x"06ad",	
												x"0690",	x"06b5",	x"06b6",	x"06be",	
												x"06ad",	x"06c8",	x"06a3",	x"06d5",	
												x"06cd",	x"06c1",	x"06e2",	x"06d4",	
												x"06eb",	x"06e0",	x"06de",	x"06e3",	
												x"06d7",	x"06e2",	x"06db",	x"06c8",	
												x"06e6",	x"06cb",	x"069e",	x"06db",	
												x"06bd",	x"06a9",	x"06d8",	x"06c8",	
												x"06ca",	x"06ae",	x"06c5",	x"06d0",	
												x"06d4",	x"06d0",	x"06e7",	x"06d3",	
												x"06d8",	x"06f0",	x"06a2",	x"06b1",	
												x"06e1",	x"06b2",	x"06f0",	x"06c7",	
												x"06e7",	x"06dd",	x"0701",	x"06f0",	
												x"06ec",	x"06c4",	x"06f6",	x"06d4",	
												x"06e3",	x"06de",	x"06ac",	x"06d2",	
												x"3030",	x"2135",	x"067a",	x"069f",	
												x"06a3",	x"0673",	x"0682",	x"0690",	
												x"06b5",	x"068c",	x"06ba",	x"069a",	
												x"06ab",	x"06c0",	x"06a8",	x"06ae",	
												x"0685",	x"06a6",	x"06bd",	x"0699",	
												x"06d9",	x"06b9",	x"06d5",	x"06da",	
												x"06dc",	x"06db",	x"06ae",	x"06c1",	
												x"06c8",	x"06cb",	x"06db",	x"06bb",	
												x"069f",	x"06c3",	x"06d9",	x"0693",	
												x"06ef",	x"06dd",	x"06d7",	x"06e6",	
												x"06d2",	x"06db",	x"06d7",	x"06c0",	
												x"06da",	x"06d0",	x"06e8",	x"06cf",	
												x"06ab",	x"06c3",	x"06ee",	x"06bc",	
												x"0700",	x"06ef",	x"06e6",	x"06de",	
												x"06fd",	x"06d1",	x"06fa",	x"06d3",	
												x"070a",	x"06d7",	x"0701",	x"06d9",	
												x"0698",	x"06eb",	x"0004",	x"000a",	
												x"0945",	x"72f3",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"2136",	
												x"06b0",	x"06ac",	x"06c1",	x"0690",	
												x"06c0",	x"06ac",	x"06c9",	x"06b5",	
												x"06cf",	x"06ba",	x"06bc",	x"06c8",	
												x"06c0",	x"06b5",	x"06ba",	x"06b6",	
												x"06df",	x"06cd",	x"06ec",	x"06db",	
												x"06f1",	x"0701",	x"0700",	x"070c",	
												x"06eb",	x"06dc",	x"06f5",	x"06d8",	
												x"06eb",	x"06f1",	x"06d7",	x"06fc",	
												x"06ff",	x"06d3",	x"0708",	x"0714",	
												x"0700",	x"06ff",	x"06e9",	x"070f",	
												x"0706",	x"0709",	x"070b",	x"0708",	
												x"0716",	x"071a",	x"0705",	x"0708",	
												x"0739",	x"06ed",	x"0708",	x"0728",	
												x"072b",	x"0703",	x"0721",	x"0718",	
												x"0721",	x"070f",	x"0728",	x"0717",	
												x"072b",	x"071f",	x"06b9",	x"071a",	
												x"5030",	x"2136",	x"06d8",	x"06bc",	
												x"06e8",	x"06da",	x"06df",	x"06c6",	
												x"06ee",	x"06d0",	x"06f2",	x"06d9",	
												x"0718",	x"06dd",	x"0701",	x"070c",	
												x"0708",	x"0702",	x"0729",	x"06fe",	
												x"072c",	x"0705",	x"0729",	x"071f",	
												x"073e",	x"0726",	x"0717",	x"070a",	
												x"072a",	x"0729",	x"0726",	x"0714",	
												x"0715",	x"070d",	x"072a",	x"070a",	
												x"0730",	x"0728",	x"072c",	x"072e",	
												x"0755",	x"0712",	x"074d",	x"072f",	
												x"074c",	x"0728",	x"074f",	x"0719",	
												x"0733",	x"0727",	x"075b",	x"0722",	
												x"0765",	x"0733",	x"077b",	x"0741",	
												x"0776",	x"0741",	x"077f",	x"074d",	
												x"0753",	x"074a",	x"0757",	x"0731",	
												x"06e9",	x"073a",	x"6030",	x"2136",	
												x"06f8",	x"06d3",	x"06eb",	x"06f9",	
												x"06f2",	x"06cf",	x"0718",	x"06f7",	
												x"071c",	x"0715",	x"0723",	x"071c",	
												x"071a",	x"0717",	x"071b",	x"06f0",	
												x"0734",	x"0703",	x"073e",	x"071c",	
												x"0745",	x"0737",	x"0762",	x"0755",	
												x"075c",	x"0760",	x"0755",	x"0742",	
												x"0750",	x"0737",	x"0734",	x"073e",	
												x"0757",	x"0723",	x"0798",	x"0755",	
												x"0761",	x"0757",	x"075d",	x"075d",	
												x"0756",	x"075b",	x"0780",	x"0735",	
												x"0761",	x"074b",	x"075f",	x"074e",	
												x"0787",	x"074d",	x"07b2",	x"0760",	
												x"078c",	x"0762",	x"079f",	x"0773",	
												x"079c",	x"0774",	x"07a7",	x"0770",	
												x"079e",	x"0775",	x"0722",	x"0775",	
												x"7030",	x"2136",	x"0772",	x"072c",	
												x"0727",	x"071c",	x"0747",	x"0710",	
												x"0773",	x"073a",	x"076d",	x"074d",	
												x"0769",	x"0754",	x"0776",	x"076b",	
												x"0773",	x"0738",	x"0792",	x"0743",	
												x"07c4",	x"0775",	x"07ad",	x"0799",	
												x"07bb",	x"07a7",	x"07b6",	x"07a8",	
												x"07f3",	x"07a1",	x"07c7",	x"07a8",	
												x"07ac",	x"0799",	x"07d4",	x"07ba",	
												x"07da",	x"07e6",	x"07d3",	x"07c7",	
												x"07d0",	x"07d5",	x"07e1",	x"07d7",	
												x"07c5",	x"07d3",	x"07dd",	x"07ca",	
												x"07de",	x"07d0",	x"07f9",	x"07d9",	
												x"07e4",	x"07e8",	x"080a",	x"07ea",	
												x"0816",	x"07ee",	x"080f",	x"07f1",	
												x"0824",	x"07f4",	x"080e",	x"07f5",	
												x"06dd",	x"07fd",	x"0004",	x"000a",	
												x"4472",	x"a446",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"3137",	
												x"0705",	x"06fb",	x"06fc",	x"0710",	
												x"06d9",	x"06f2",	x"06fc",	x"06fa",	
												x"072b",	x"071d",	x"0723",	x"070a",	
												x"0718",	x"0710",	x"0705",	x"0717",	
												x"0738",	x"073e",	x"0753",	x"076c",	
												x"071b",	x"0751",	x"0743",	x"0743",	
												x"073f",	x"0757",	x"0721",	x"074a",	
												x"0723",	x"0732",	x"06d3",	x"071a",	
												x"0726",	x"0718",	x"0738",	x"0739",	
												x"072d",	x"0744",	x"072c",	x"0745",	
												x"0747",	x"0734",	x"0731",	x"0739",	
												x"071c",	x"072d",	x"06f7",	x"072b",	
												x"0723",	x"06fd",	x"0755",	x"0753",	
												x"075e",	x"0753",	x"0750",	x"077a",	
												x"0734",	x"075c",	x"0742",	x"0744",	
												x"0719",	x"071b",	x"06b0",	x"071a",	
												x"1030",	x"3137",	x"06a9",	x"06e0",	
												x"06fc",	x"06d8",	x"06c2",	x"06e4",	
												x"06cb",	x"06db",	x"0700",	x"06ea",	
												x"0706",	x"0717",	x"070c",	x"0715",	
												x"06ce",	x"0712",	x"0719",	x"06f8",	
												x"073e",	x"0724",	x"071d",	x"073b",	
												x"075a",	x"0756",	x"0708",	x"073d",	
												x"0733",	x"0729",	x"072c",	x"0711",	
												x"06da",	x"0716",	x"070f",	x"06f1",	
												x"0715",	x"0722",	x"0738",	x"0722",	
												x"073c",	x"074f",	x"072f",	x"072b",	
												x"0712",	x"0721",	x"06f9",	x"0712",	
												x"06fd",	x"0708",	x"071c",	x"06fd",	
												x"0725",	x"0711",	x"0738",	x"0735",	
												x"0748",	x"0745",	x"0737",	x"0742",	
												x"071f",	x"073c",	x"073c",	x"0725",	
												x"06da",	x"0722",	x"2030",	x"3137",	
												x"06b3",	x"0718",	x"06c1",	x"06d2",	
												x"06bc",	x"06ff",	x"06d2",	x"06e5",	
												x"071a",	x"06f3",	x"06de",	x"06f8",	
												x"06f2",	x"0703",	x"06bc",	x"070f",	
												x"0704",	x"06fb",	x"0711",	x"0734",	
												x"072d",	x"072c",	x"06f8",	x"072c",	
												x"06fb",	x"0714",	x"06f6",	x"0718",	
												x"06fb",	x"06f3",	x"06d0",	x"06fe",	
												x"0708",	x"06f9",	x"0710",	x"071c",	
												x"0721",	x"072b",	x"0711",	x"0710",	
												x"072b",	x"0718",	x"071b",	x"0716",	
												x"070d",	x"0708",	x"06dd",	x"06fa",	
												x"071d",	x"06ee",	x"0716",	x"070c",	
												x"071f",	x"0726",	x"071b",	x"071e",	
												x"071b",	x"0706",	x"0724",	x"0717",	
												x"072c",	x"06fb",	x"06bb",	x"06f8",	
												x"3030",	x"3137",	x"06c0",	x"06c8",	
												x"06a1",	x"06cf",	x"06b4",	x"06ba",	
												x"06ac",	x"06c9",	x"06c9",	x"06ae",	
												x"06ed",	x"06d9",	x"06dd",	x"06cc",	
												x"06c1",	x"06e6",	x"06e8",	x"06d6",	
												x"06fd",	x"06ef",	x"0719",	x"0704",	
												x"0706",	x"0706",	x"0707",	x"06e2",	
												x"0717",	x"06ff",	x"06f4",	x"0703",	
												x"0697",	x"06ea",	x"06f7",	x"06c2",	
												x"070e",	x"06fe",	x"071c",	x"06f9",	
												x"0711",	x"0720",	x"06fb",	x"070a",	
												x"070c",	x"06f4",	x"0705",	x"06f3",	
												x"06f5",	x"06ff",	x"071c",	x"06fc",	
												x"0717",	x"0717",	x"071a",	x"070d",	
												x"072f",	x"071b",	x"071c",	x"0722",	
												x"0716",	x"0715",	x"071d",	x"0705",	
												x"06c9",	x"070b",	x"0004",	x"000a",	
												x"2414",	x"d154",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"3138",	
												x"06d4",	x"06f7",	x"06d8",	x"06c7",	
												x"06d6",	x"06cb",	x"06e2",	x"06da",	
												x"06ed",	x"06d2",	x"071d",	x"06dd",	
												x"06f5",	x"070f",	x"06ff",	x"0704",	
												x"0716",	x"070f",	x"0746",	x"072d",	
												x"071e",	x"0725",	x"0726",	x"0738",	
												x"072f",	x"070e",	x"0728",	x"073d",	
												x"0711",	x"0709",	x"0709",	x"071c",	
												x"0730",	x"06f9",	x"072c",	x"073e",	
												x"074c",	x"072c",	x"0756",	x"0753",	
												x"0724",	x"073a",	x"0742",	x"0734",	
												x"0745",	x"0739",	x"072d",	x"073b",	
												x"0741",	x"072f",	x"0763",	x"0742",	
												x"0773",	x"0762",	x"0777",	x"0773",	
												x"0766",	x"0763",	x"076b",	x"0762",	
												x"075a",	x"0761",	x"070f",	x"0752",	
												x"5030",	x"3138",	x"0721",	x"070a",	
												x"072a",	x"06f5",	x"072b",	x"0715",	
												x"0732",	x"0731",	x"074c",	x"0718",	
												x"0746",	x"0731",	x"0735",	x"073e",	
												x"073c",	x"072e",	x"0764",	x"0740",	
												x"0763",	x"0752",	x"0763",	x"0753",	
												x"0777",	x"0763",	x"0763",	x"0759",	
												x"077b",	x"075e",	x"075e",	x"074c",	
												x"0741",	x"074a",	x"0771",	x"0728",	
												x"077c",	x"0773",	x"0776",	x"0754",	
												x"0789",	x"0771",	x"076e",	x"075f",	
												x"0775",	x"0762",	x"078d",	x"0737",	
												x"076c",	x"0747",	x"07a7",	x"073b",	
												x"07af",	x"076a",	x"07a7",	x"0779",	
												x"07ae",	x"077e",	x"079b",	x"077f",	
												x"07a3",	x"0767",	x"0792",	x"076f",	
												x"0726",	x"0749",	x"6030",	x"3138",	
												x"0746",	x"06f8",	x"0750",	x"0703",	
												x"0704",	x"0728",	x"075b",	x"070c",	
												x"0766",	x"073e",	x"075d",	x"073e",	
												x"0750",	x"0759",	x"0738",	x"0742",	
												x"076c",	x"0735",	x"079d",	x"0749",	
												x"079f",	x"076a",	x"0793",	x"0777",	
												x"078e",	x"078f",	x"0787",	x"076a",	
												x"0788",	x"0757",	x"0768",	x"0760",	
												x"07a8",	x"0772",	x"07b5",	x"07a1",	
												x"07a6",	x"0791",	x"07c7",	x"07ad",	
												x"07a2",	x"0796",	x"07ab",	x"0794",	
												x"07a8",	x"0792",	x"07ab",	x"079d",	
												x"07d7",	x"0793",	x"07e0",	x"07b7",	
												x"07cf",	x"07a4",	x"07e5",	x"07ac",	
												x"07cb",	x"0793",	x"07c3",	x"078a",	
												x"07db",	x"0794",	x"0775",	x"079e",	
												x"7030",	x"3138",	x"0795",	x"076a",	
												x"079d",	x"0782",	x"0797",	x"0796",	
												x"0785",	x"0771",	x"0767",	x"0752",	
												x"07b1",	x"0763",	x"07b2",	x"07b4",	
												x"07a2",	x"07be",	x"0803",	x"0792",	
												x"0800",	x"07df",	x"0810",	x"07f5",	
												x"0816",	x"07e9",	x"080a",	x"07eb",	
												x"07f4",	x"07f6",	x"0806",	x"07d6",	
												x"07df",	x"07ec",	x"0802",	x"07e8",	
												x"0814",	x"080e",	x"081e",	x"0800",	
												x"0840",	x"080d",	x"081f",	x"0829",	
												x"081d",	x"081b",	x"0818",	x"07e6",	
												x"0832",	x"082c",	x"0839",	x"0827",	
												x"0841",	x"082d",	x"0845",	x"0826",	
												x"0878",	x"0844",	x"0881",	x"0820",	
												x"0872",	x"0838",	x"0846",	x"083d",	
												x"0660",	x"0828",	x"0004",	x"000a",	
												x"62a2",	x"0184",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"0139",	
												x"065f",	x"0690",	x"0664",	x"0658",	
												x"064a",	x"0668",	x"0648",	x"0644",	
												x"0653",	x"0642",	x"0643",	x"063a",	
												x"0645",	x"063e",	x"0634",	x"0647",	
												x"066d",	x"062b",	x"0696",	x"064e",	
												x"0699",	x"067a",	x"0691",	x"06b6",	
												x"0668",	x"0671",	x"0675",	x"067d",	
												x"0669",	x"065f",	x"0645",	x"0676",	
												x"0666",	x"0651",	x"0692",	x"0675",	
												x"066b",	x"0688",	x"0689",	x"0697",	
												x"0695",	x"0674",	x"068a",	x"0688",	
												x"0667",	x"068d",	x"0655",	x"0685",	
												x"0686",	x"0663",	x"0678",	x"0688",	
												x"0679",	x"067f",	x"0689",	x"0675",	
												x"0687",	x"0682",	x"06cb",	x"0687",	
												x"067e",	x"068e",	x"062d",	x"0670",	
												x"1031",	x"0139",	x"0633",	x"066f",	
												x"065a",	x"0653",	x"0633",	x"0659",	
												x"0639",	x"0645",	x"0628",	x"063b",	
												x"0630",	x"0621",	x"061b",	x"0619",	
												x"062d",	x"0628",	x"0660",	x"064a",	
												x"067b",	x"0658",	x"067f",	x"066a",	
												x"0664",	x"0682",	x"0669",	x"067f",	
												x"0667",	x"067d",	x"0667",	x"0670",	
												x"0630",	x"066e",	x"068b",	x"063d",	
												x"0652",	x"0680",	x"0671",	x"066c",	
												x"0685",	x"0689",	x"067d",	x"068c",	
												x"0672",	x"067c",	x"066b",	x"0663",	
												x"0658",	x"0671",	x"0656",	x"0667",	
												x"0694",	x"0694",	x"0694",	x"06a1",	
												x"068d",	x"0697",	x"0689",	x"0686",	
												x"0694",	x"0698",	x"0688",	x"068d",	
												x"063c",	x"0687",	x"2031",	x"0139",	
												x"0635",	x"0632",	x"0665",	x"0641",	
												x"0629",	x"064c",	x"0626",	x"0623",	
												x"061a",	x"0638",	x"0646",	x"064a",	
												x"0649",	x"0650",	x"0617",	x"0659",	
												x"0636",	x"064b",	x"0662",	x"0662",	
												x"0681",	x"0673",	x"066c",	x"0672",	
												x"064f",	x"0673",	x"0649",	x"0672",	
												x"0654",	x"064c",	x"0632",	x"0659",	
												x"0654",	x"0663",	x"0663",	x"0663",	
												x"065d",	x"065d",	x"0661",	x"0681",	
												x"066c",	x"0662",	x"0668",	x"065e",	
												x"0661",	x"065b",	x"0653",	x"065b",	
												x"0672",	x"065c",	x"067c",	x"0660",	
												x"0679",	x"066d",	x"0678",	x"0694",	
												x"065e",	x"0681",	x"0675",	x"067d",	
												x"067d",	x"066f",	x"0622",	x"0675",	
												x"3031",	x"0139",	x"0642",	x"063e",	
												x"063c",	x"061d",	x"0628",	x"061b",	
												x"0625",	x"061e",	x"061e",	x"060c",	
												x"061f",	x"0619",	x"0632",	x"061a",	
												x"0621",	x"0632",	x"065e",	x"0627",	
												x"0662",	x"0651",	x"065d",	x"064f",	
												x"065c",	x"0670",	x"0642",	x"0645",	
												x"066b",	x"0649",	x"0657",	x"0657",	
												x"0651",	x"0654",	x"0654",	x"064f",	
												x"0671",	x"064e",	x"0669",	x"0655",	
												x"0675",	x"066d",	x"0683",	x"064a",	
												x"068a",	x"0670",	x"067a",	x"0677",	
												x"065f",	x"0651",	x"066e",	x"064c",	
												x"0683",	x"064c",	x"0692",	x"0669",	
												x"0693",	x"067e",	x"06a1",	x"066d",	
												x"06a7",	x"0669",	x"068d",	x"066f",	
												x"062b",	x"0670",	x"0004",	x"000a",	
												x"d011",	x"b970",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"013a",	
												x"0626",	x"063d",	x"0649",	x"062f",	
												x"0639",	x"064a",	x"0631",	x"0637",	
												x"0645",	x"0603",	x"0648",	x"0639",	
												x"0668",	x"063f",	x"062e",	x"063f",	
												x"0667",	x"0630",	x"067b",	x"0643",	
												x"0688",	x"0664",	x"0679",	x"0691",	
												x"0685",	x"0671",	x"0683",	x"067a",	
												x"06a1",	x"0687",	x"066a",	x"0673",	
												x"06c1",	x"066c",	x"06b7",	x"06ac",	
												x"0699",	x"069c",	x"06c3",	x"06a5",	
												x"06c3",	x"0692",	x"06bb",	x"06c1",	
												x"068f",	x"0691",	x"069c",	x"069b",	
												x"06bb",	x"068f",	x"06cf",	x"06a1",	
												x"06d6",	x"06b4",	x"06d3",	x"06cb",	
												x"06e0",	x"06c9",	x"06de",	x"06c7",	
												x"06b9",	x"06b7",	x"065b",	x"06b1",	
												x"5031",	x"013a",	x"068a",	x"066b",	
												x"0692",	x"0673",	x"067a",	x"0683",	
												x"067f",	x"067a",	x"0693",	x"0656",	
												x"0690",	x"066d",	x"06a6",	x"0679",	
												x"06a2",	x"068c",	x"06b4",	x"067e",	
												x"06c1",	x"06af",	x"06d2",	x"06bc",	
												x"06f5",	x"06ce",	x"06b6",	x"06a6",	
												x"06c8",	x"06b0",	x"06cb",	x"06af",	
												x"06bd",	x"069c",	x"06e6",	x"06a4",	
												x"06dd",	x"06a8",	x"06e5",	x"06a0",	
												x"06dd",	x"06c2",	x"06fd",	x"06c1",	
												x"06e7",	x"06c4",	x"06dc",	x"06c0",	
												x"06ca",	x"06ae",	x"06fc",	x"06ae",	
												x"06f2",	x"06c8",	x"06e3",	x"06c1",	
												x"070b",	x"06ad",	x"0704",	x"06d0",	
												x"0709",	x"06d3",	x"06e4",	x"06de",	
												x"0691",	x"06c9",	x"6031",	x"013a",	
												x"06ae",	x"0673",	x"06ac",	x"0690",	
												x"069d",	x"067f",	x"069e",	x"067a",	
												x"0693",	x"0686",	x"068a",	x"0687",	
												x"068d",	x"0677",	x"069e",	x"065a",	
												x"06e2",	x"0679",	x"06e0",	x"06be",	
												x"06df",	x"06cf",	x"06e3",	x"06e1",	
												x"06f7",	x"06d7",	x"0713",	x"06d5",	
												x"0704",	x"06c8",	x"06ea",	x"06e8",	
												x"0716",	x"06e4",	x"06fe",	x"06c4",	
												x"0711",	x"06e8",	x"0717",	x"06f9",	
												x"0717",	x"06ee",	x"072b",	x"06f5",	
												x"0742",	x"0715",	x"06f2",	x"06f5",	
												x"0735",	x"06e0",	x"072d",	x"06f4",	
												x"0749",	x"06f7",	x"072e",	x"06ff",	
												x"074a",	x"0712",	x"0738",	x"0707",	
												x"0730",	x"0705",	x"06c5",	x"06f2",	
												x"7031",	x"013a",	x"06f8",	x"06b1",	
												x"0704",	x"06ac",	x"06c2",	x"06a9",	
												x"06e3",	x"06a5",	x"06dd",	x"06a1",	
												x"071f",	x"06bc",	x"06f2",	x"06dd",	
												x"06c8",	x"06d4",	x"072f",	x"06c1",	
												x"075f",	x"0720",	x"073c",	x"072a",	
												x"074f",	x"0720",	x"074d",	x"072d",	
												x"0761",	x"071c",	x"0768",	x"0734",	
												x"071c",	x"0734",	x"0773",	x"072f",	
												x"0772",	x"0764",	x"0781",	x"074b",	
												x"0789",	x"074a",	x"0794",	x"0765",	
												x"0797",	x"0760",	x"0787",	x"077f",	
												x"076e",	x"075c",	x"079d",	x"075c",	
												x"07c6",	x"0765",	x"07a2",	x"078e",	
												x"07cd",	x"07a8",	x"07a1",	x"07af",	
												x"07cd",	x"077a",	x"079e",	x"0782",	
												x"0717",	x"0791",	x"0004",	x"000a",	
												x"1344",	x"ec12",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"113b",	
												x"074f",	x"0753",	x"074f",	x"0772",	
												x"0767",	x"0765",	x"073f",	x"077d",	
												x"071f",	x"072e",	x"0722",	x"0716",	
												x"0726",	x"0704",	x"06e0",	x"0703",	
												x"0716",	x"06df",	x"06f1",	x"0723",	
												x"072b",	x"0728",	x"0739",	x"073b",	
												x"073a",	x"074b",	x"0770",	x"0765",	
												x"0725",	x"0764",	x"071e",	x"077a",	
												x"074f",	x"071f",	x"0738",	x"0784",	
												x"073d",	x"073c",	x"073d",	x"075d",	
												x"073e",	x"074f",	x"0745",	x"0750",	
												x"076f",	x"0746",	x"06e2",	x"0761",	
												x"0739",	x"070d",	x"0744",	x"0738",	
												x"0758",	x"0741",	x"0761",	x"0755",	
												x"073e",	x"072e",	x"0758",	x"073c",	
												x"0748",	x"073a",	x"072d",	x"0754",	
												x"1031",	x"113b",	x"073e",	x"0739",	
												x"074b",	x"0759",	x"073c",	x"0752",	
												x"0718",	x"074f",	x"072e",	x"070b",	
												x"06e9",	x"0708",	x"06fe",	x"06da",	
												x"06cb",	x"06f1",	x"06e5",	x"06d6",	
												x"0702",	x"06ee",	x"0709",	x"06f8",	
												x"0717",	x"0704",	x"074f",	x"0748",	
												x"0719",	x"0741",	x"0744",	x"074d",	
												x"072b",	x"0759",	x"0754",	x"0726",	
												x"0767",	x"0760",	x"0748",	x"074d",	
												x"0737",	x"0752",	x"0736",	x"0757",	
												x"0759",	x"074c",	x"0756",	x"0750",	
												x"070e",	x"0756",	x"0731",	x"0714",	
												x"0740",	x"073e",	x"0738",	x"0741",	
												x"0749",	x"0750",	x"073d",	x"0747",	
												x"0772",	x"076a",	x"0777",	x"075d",	
												x"071d",	x"0748",	x"2031",	x"113b",	
												x"0741",	x"072c",	x"071f",	x"0709",	
												x"072e",	x"0716",	x"071c",	x"0737",	
												x"0703",	x"0722",	x"06fe",	x"070f",	
												x"06f6",	x"0704",	x"06ca",	x"06f0",	
												x"06e3",	x"06f4",	x"06f9",	x"0703",	
												x"06e9",	x"06ef",	x"06f2",	x"06fc",	
												x"0729",	x"0717",	x"071d",	x"0739",	
												x"071f",	x"071a",	x"06f9",	x"0719",	
												x"0722",	x"06f8",	x"074f",	x"0721",	
												x"072c",	x"0736",	x"0724",	x"072c",	
												x"0740",	x"071c",	x"074b",	x"072b",	
												x"0727",	x"072a",	x"06ef",	x"0719",	
												x"0733",	x"0704",	x"0723",	x"0729",	
												x"0722",	x"072f",	x"0741",	x"0740",	
												x"0748",	x"071c",	x"074b",	x"0745",	
												x"0742",	x"0746",	x"06f1",	x"073b",	
												x"3031",	x"113b",	x"0715",	x"06eb",	
												x"0702",	x"06ee",	x"0700",	x"06e7",	
												x"06ff",	x"0712",	x"06e4",	x"06f4",	
												x"06f8",	x"06d2",	x"06db",	x"06df",	
												x"06e3",	x"06c8",	x"06ed",	x"06d2",	
												x"06ed",	x"06e7",	x"0706",	x"06c6",	
												x"0732",	x"0708",	x"0735",	x"0716",	
												x"0745",	x"072b",	x"0718",	x"072e",	
												x"071a",	x"070e",	x"0747",	x"0707",	
												x"071c",	x"072b",	x"076c",	x"0725",	
												x"0743",	x"073d",	x"0737",	x"0737",	
												x"073f",	x"0730",	x"0753",	x"073c",	
												x"0725",	x"072a",	x"075d",	x"0715",	
												x"0751",	x"0734",	x"0746",	x"0722",	
												x"0750",	x"0736",	x"0763",	x"0734",	
												x"0762",	x"072f",	x"075c",	x"0723",	
												x"0717",	x"072d",	x"0004",	x"000a",	
												x"34e1",	x"5d43",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"113c",	
												x"0738",	x"06fb",	x"0746",	x"0720",	
												x"0728",	x"0724",	x"072d",	x"0716",	
												x"0727",	x"06ec",	x"071f",	x"0708",	
												x"070a",	x"06f4",	x"06d7",	x"06cc",	
												x"070c",	x"06e2",	x"0716",	x"06d6",	
												x"072a",	x"0715",	x"0769",	x"072a",	
												x"0755",	x"0714",	x"076b",	x"0747",	
												x"0751",	x"074c",	x"074f",	x"073c",	
												x"076f",	x"0749",	x"0792",	x"0768",	
												x"0798",	x"077f",	x"0769",	x"0751",	
												x"0785",	x"0770",	x"0781",	x"076a",	
												x"077d",	x"0771",	x"076c",	x"0764",	
												x"07a5",	x"075b",	x"07b1",	x"0776",	
												x"0782",	x"0764",	x"0781",	x"0778",	
												x"079f",	x"0765",	x"07bc",	x"0783",	
												x"07a8",	x"078a",	x"0748",	x"077a",	
												x"5031",	x"113c",	x"0765",	x"074d",	
												x"0772",	x"074a",	x"075e",	x"075a",	
												x"078f",	x"0765",	x"074f",	x"0737",	
												x"073a",	x"0756",	x"0742",	x"0744",	
												x"073a",	x"0734",	x"0754",	x"0709",	
												x"0761",	x"0750",	x"0782",	x"075b",	
												x"0791",	x"0766",	x"079d",	x"0793",	
												x"0799",	x"074f",	x"07a0",	x"0784",	
												x"078b",	x"076c",	x"079f",	x"0753",	
												x"07af",	x"0785",	x"07a5",	x"0768",	
												x"07a2",	x"0775",	x"07b6",	x"078b",	
												x"07d1",	x"078c",	x"07cf",	x"078a",	
												x"07b7",	x"078e",	x"07c3",	x"0765",	
												x"07cc",	x"07a9",	x"07cd",	x"0792",	
												x"07d0",	x"0786",	x"07d0",	x"0795",	
												x"07fc",	x"078e",	x"07c2",	x"079e",	
												x"0751",	x"0790",	x"6031",	x"113c",	
												x"076d",	x"074d",	x"077b",	x"074e",	
												x"0781",	x"0753",	x"0771",	x"0768",	
												x"077e",	x"074b",	x"077c",	x"0748",	
												x"0769",	x"0752",	x"073b",	x"0714",	
												x"078a",	x"071d",	x"07b3",	x"0751",	
												x"079b",	x"0756",	x"07d4",	x"0793",	
												x"07bb",	x"07a1",	x"07be",	x"0792",	
												x"07d4",	x"0795",	x"07bf",	x"077e",	
												x"07db",	x"077e",	x"07f2",	x"07ad",	
												x"07e0",	x"07b1",	x"07dc",	x"07c5",	
												x"07f5",	x"07b1",	x"07fc",	x"07c0",	
												x"07e0",	x"07cc",	x"07cd",	x"07b4",	
												x"07f7",	x"07a6",	x"07f8",	x"07de",	
												x"080a",	x"07c0",	x"07fd",	x"07c1",	
												x"0833",	x"07bf",	x"080c",	x"07bc",	
												x"0819",	x"07ac",	x"079a",	x"07c7",	
												x"7031",	x"113c",	x"07bb",	x"078a",	
												x"07bb",	x"079b",	x"07d0",	x"0792",	
												x"07d8",	x"0799",	x"07bd",	x"07a2",	
												x"07ca",	x"07a0",	x"07a2",	x"07a5",	
												x"079a",	x"079c",	x"07e2",	x"0775",	
												x"07cc",	x"078e",	x"0813",	x"07b1",	
												x"0817",	x"07b2",	x"082b",	x"07e5",	
												x"0837",	x"0815",	x"0838",	x"07f5",	
												x"0840",	x"0801",	x"086a",	x"07cb",	
												x"0863",	x"082a",	x"0872",	x"082f",	
												x"0876",	x"0829",	x"0857",	x"083b",	
												x"0862",	x"0836",	x"0889",	x"0848",	
												x"0844",	x"082f",	x"0858",	x"0841",	
												x"086e",	x"085b",	x"086a",	x"0858",	
												x"085e",	x"085b",	x"089c",	x"0850",	
												x"08a2",	x"086c",	x"088b",	x"0877",	
												x"06c7",	x"0857",	x"0004",	x"000a",	
												x"7a0e",	x"8ed6",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"213d",	
												x"06e2",	x"06dd",	x"06e3",	x"0707",	
												x"06f2",	x"06e9",	x"070a",	x"06e5",	
												x"06a5",	x"06e9",	x"06b7",	x"06b1",	
												x"06a8",	x"06c5",	x"067e",	x"0698",	
												x"069a",	x"0684",	x"06b3",	x"06c8",	
												x"06eb",	x"06e3",	x"0703",	x"070d",	
												x"06fa",	x"0715",	x"0702",	x"0701",	
												x"06ea",	x"070a",	x"06ab",	x"06f7",	
												x"06e1",	x"06d0",	x"06e7",	x"06f5",	
												x"06f8",	x"06f5",	x"06ee",	x"0706",	
												x"06f4",	x"06f9",	x"06df",	x"06f3",	
												x"0705",	x"06e5",	x"06b7",	x"06db",	
												x"06e6",	x"06da",	x"06ee",	x"0708",	
												x"06f3",	x"06e4",	x"06f8",	x"06ef",	
												x"0710",	x"06ea",	x"072b",	x"06f6",	
												x"071a",	x"0716",	x"06be",	x"0716",	
												x"1031",	x"213d",	x"06c6",	x"06d2",	
												x"06d7",	x"06da",	x"06ce",	x"06cc",	
												x"06cb",	x"06dd",	x"06c1",	x"06c6",	
												x"06bb",	x"06a8",	x"0678",	x"067d",	
												x"0650",	x"0658",	x"0675",	x"0673",	
												x"06bd",	x"0667",	x"06be",	x"06a6",	
												x"06d6",	x"06b4",	x"06c7",	x"06d6",	
												x"070e",	x"06de",	x"06c5",	x"0703",	
												x"0694",	x"06dc",	x"06d7",	x"069f",	
												x"06d6",	x"06e5",	x"06de",	x"06de",	
												x"06d7",	x"06f1",	x"06e7",	x"06e5",	
												x"06e7",	x"06f9",	x"06eb",	x"06e5",	
												x"06b6",	x"06e3",	x"06e7",	x"06df",	
												x"06e2",	x"06d9",	x"06e8",	x"06d9",	
												x"06f8",	x"06e6",	x"070a",	x"06e1",	
												x"0727",	x"06ee",	x"070a",	x"072b",	
												x"06ac",	x"06fa",	x"2031",	x"213d",	
												x"06a9",	x"06e0",	x"06b0",	x"06bc",	
												x"06b7",	x"06c6",	x"06a3",	x"06d8",	
												x"0693",	x"06bb",	x"0697",	x"0693",	
												x"0692",	x"0681",	x"063b",	x"0688",	
												x"0689",	x"066d",	x"0681",	x"06a0",	
												x"06c4",	x"06a3",	x"06ce",	x"06d5",	
												x"06ec",	x"06d2",	x"06cc",	x"06d2",	
												x"06bf",	x"06d7",	x"06bc",	x"06bf",	
												x"06cc",	x"06bd",	x"06fd",	x"06d2",	
												x"06d1",	x"06d7",	x"06d3",	x"06d1",	
												x"06cd",	x"06b2",	x"06df",	x"06d1",	
												x"06ed",	x"06e9",	x"06b9",	x"06d6",	
												x"06d8",	x"06c4",	x"06bf",	x"06ca",	
												x"06dc",	x"06c5",	x"06e9",	x"06f4",	
												x"06e8",	x"06cf",	x"070e",	x"06df",	
												x"06fc",	x"06ed",	x"069c",	x"06f4",	
												x"3031",	x"213d",	x"06a3",	x"0691",	
												x"06ad",	x"0693",	x"06a9",	x"06ae",	
												x"06b7",	x"069b",	x"06af",	x"0690",	
												x"0691",	x"0697",	x"066c",	x"068a",	
												x"065f",	x"067e",	x"069a",	x"0668",	
												x"06bd",	x"068c",	x"06bc",	x"06c4",	
												x"06e4",	x"06bd",	x"06d0",	x"06ba",	
												x"06d1",	x"06d0",	x"06e1",	x"06b3",	
												x"06b5",	x"06b9",	x"06d7",	x"06a2",	
												x"06f5",	x"06bc",	x"06e0",	x"06d4",	
												x"06de",	x"06ce",	x"06ed",	x"06c3",	
												x"06dc",	x"06dc",	x"06db",	x"06db",	
												x"06ca",	x"06c2",	x"0704",	x"06c3",	
												x"06cb",	x"06d5",	x"06e2",	x"06c2",	
												x"06f1",	x"06ca",	x"06ff",	x"06d6",	
												x"0721",	x"06d9",	x"071c",	x"0704",	
												x"06a1",	x"06eb",	x"0004",	x"000a",	
												x"070f",	x"6f73",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"213e",	
												x"06c3",	x"06ad",	x"06d7",	x"06be",	
												x"06e1",	x"06bb",	x"06c9",	x"06c1",	
												x"06b6",	x"06bf",	x"06a7",	x"06aa",	
												x"06a2",	x"068d",	x"0694",	x"06b6",	
												x"06d6",	x"0665",	x"06e5",	x"06be",	
												x"06ef",	x"06f1",	x"0711",	x"06fa",	
												x"0700",	x"06ed",	x"070f",	x"0701",	
												x"0704",	x"0703",	x"06e3",	x"06fc",	
												x"06fb",	x"06d6",	x"072c",	x"0716",	
												x"074e",	x"0710",	x"072b",	x"0712",	
												x"0722",	x"071c",	x"072c",	x"0706",	
												x"072f",	x"0725",	x"0713",	x"0726",	
												x"0726",	x"06fc",	x"0733",	x"070e",	
												x"073c",	x"070d",	x"0748",	x"071e",	
												x"0765",	x"070d",	x"0768",	x"0732",	
												x"0774",	x"0740",	x"06c3",	x"073b",	
												x"5031",	x"213e",	x"070e",	x"06d0",	
												x"070f",	x"0708",	x"0715",	x"06d8",	
												x"0714",	x"070a",	x"0719",	x"06ea",	
												x"06fa",	x"06cf",	x"06fd",	x"06ce",	
												x"06fe",	x"06f0",	x"0706",	x"06bb",	
												x"074f",	x"06fa",	x"073a",	x"0711",	
												x"0753",	x"0731",	x"072d",	x"070a",	
												x"072a",	x"0725",	x"0742",	x"0715",	
												x"071c",	x"070f",	x"0740",	x"0706",	
												x"073e",	x"073a",	x"074e",	x"0705",	
												x"075c",	x"0731",	x"0774",	x"0732",	
												x"0778",	x"0745",	x"0766",	x"0747",	
												x"0738",	x"072d",	x"076a",	x"072d",	
												x"0762",	x"074e",	x"075c",	x"071f",	
												x"0796",	x"072a",	x"0796",	x"0737",	
												x"078c",	x"0766",	x"0776",	x"0749",	
												x"0700",	x"0748",	x"6031",	x"213e",	
												x"0738",	x"06f9",	x"0719",	x"06f8",	
												x"0728",	x"06dc",	x"0713",	x"06e5",	
												x"0706",	x"06df",	x"0709",	x"06df",	
												x"0705",	x"06f3",	x"0708",	x"06dc",	
												x"0725",	x"06b8",	x"0734",	x"06fc",	
												x"075d",	x"0707",	x"0781",	x"0734",	
												x"077e",	x"0753",	x"0773",	x"0750",	
												x"0779",	x"072b",	x"074f",	x"0744",	
												x"0792",	x"0743",	x"0789",	x"0780",	
												x"0782",	x"0776",	x"079f",	x"0766",	
												x"0797",	x"0763",	x"07a3",	x"076f",	
												x"0793",	x"0770",	x"0789",	x"0760",	
												x"0780",	x"0758",	x"07b1",	x"0762",	
												x"07a1",	x"0761",	x"07c3",	x"0757",	
												x"07e3",	x"0767",	x"07e4",	x"0779",	
												x"07e1",	x"077e",	x"0755",	x"077e",	
												x"7031",	x"213e",	x"0790",	x"072a",	
												x"0760",	x"0754",	x"0772",	x"0738",	
												x"076b",	x"0759",	x"0745",	x"0743",	
												x"074a",	x"074b",	x"0761",	x"0736",	
												x"0734",	x"0711",	x"0799",	x"06e8",	
												x"07a4",	x"071d",	x"07bf",	x"075b",	
												x"07d7",	x"07a9",	x"07f8",	x"0790",	
												x"07f1",	x"079b",	x"07f7",	x"07ab",	
												x"07be",	x"07b3",	x"07f2",	x"07b4",	
												x"07e2",	x"07b1",	x"07ff",	x"07bc",	
												x"081c",	x"07f2",	x"0804",	x"07b7",	
												x"0801",	x"07e8",	x"082d",	x"07dd",	
												x"07d4",	x"07e6",	x"0815",	x"07c2",	
												x"07f0",	x"07e7",	x"07ee",	x"07eb",	
												x"083d",	x"07f1",	x"082b",	x"07ea",	
												x"0830",	x"0806",	x"0826",	x"07fb",	
												x"071d",	x"0810",	x"0004",	x"000a",	
												x"4f0d",	x"a3e8",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"313f",	
												x"0732",	x"072b",	x"073e",	x"0743",	
												x"0735",	x"0736",	x"0738",	x"0739",	
												x"0718",	x"0714",	x"0720",	x"070a",	
												x"06fc",	x"0701",	x"06ac",	x"06d8",	
												x"06de",	x"06d5",	x"06e2",	x"06ed",	
												x"06df",	x"06ef",	x"0719",	x"074c",	
												x"0734",	x"0723",	x"0744",	x"073d",	
												x"0720",	x"0745",	x"06f7",	x"0725",	
												x"0717",	x"0712",	x"073d",	x"0746",	
												x"072d",	x"0757",	x"071b",	x"0752",	
												x"070f",	x"06fa",	x"0733",	x"06ff",	
												x"0742",	x"0721",	x"0701",	x"0736",	
												x"071a",	x"0726",	x"0728",	x"0732",	
												x"0725",	x"073a",	x"0724",	x"072d",	
												x"074d",	x"0724",	x"0756",	x"071f",	
												x"0748",	x"072f",	x"06ec",	x"0736",	
												x"1031",	x"313f",	x"0725",	x"071f",	
												x"0723",	x"074a",	x"0706",	x"0719",	
												x"071e",	x"0714",	x"06ea",	x"0716",	
												x"06ea",	x"06f3",	x"06bb",	x"06ee",	
												x"06b0",	x"06c4",	x"06d0",	x"06a9",	
												x"0703",	x"06bb",	x"06ff",	x"0713",	
												x"070c",	x"0717",	x"0711",	x"0716",	
												x"072b",	x"0739",	x"0727",	x"0728",	
												x"06c8",	x"0729",	x"0714",	x"0708",	
												x"0727",	x"0743",	x"0718",	x"0726",	
												x"0758",	x"073c",	x"0719",	x"0740",	
												x"071a",	x"073b",	x"0730",	x"0712",	
												x"0702",	x"0739",	x"072d",	x"0718",	
												x"073c",	x"072b",	x"0720",	x"072e",	
												x"0720",	x"074a",	x"072d",	x"0709",	
												x"073e",	x"072d",	x"0749",	x"072d",	
												x"06de",	x"0723",	x"2031",	x"313f",	
												x"06f7",	x"070f",	x"06e6",	x"0719",	
												x"0703",	x"070f",	x"06f2",	x"071e",	
												x"06df",	x"06ef",	x"06e9",	x"06db",	
												x"06ae",	x"06c5",	x"0662",	x"06ae",	
												x"06db",	x"069d",	x"06d1",	x"06d8",	
												x"06e1",	x"06f4",	x"06df",	x"06f4",	
												x"0704",	x"06f0",	x"0708",	x"0711",	
												x"0712",	x"06f9",	x"06e6",	x"070d",	
												x"0737",	x"0702",	x"06fe",	x"0739",	
												x"071d",	x"0708",	x"071a",	x"06f2",	
												x"0721",	x"0712",	x"0725",	x"0723",	
												x"0708",	x"0707",	x"0709",	x"0718",	
												x"0733",	x"06f8",	x"0701",	x"070a",	
												x"0719",	x"0715",	x"0715",	x"0729",	
												x"0711",	x"06ed",	x"0740",	x"0715",	
												x"0740",	x"0713",	x"06b3",	x"06fb",	
												x"3031",	x"313f",	x"06dc",	x"06bb",	
												x"06e8",	x"06d8",	x"070e",	x"06f1",	
												x"0706",	x"06fd",	x"06cf",	x"06c1",	
												x"06ea",	x"06bd",	x"06a7",	x"0699",	
												x"06b2",	x"06b9",	x"06c3",	x"06ad",	
												x"06c4",	x"068b",	x"06ec",	x"06c7",	
												x"0711",	x"06d3",	x"0715",	x"06f7",	
												x"0718",	x"0703",	x"0723",	x"06f6",	
												x"06db",	x"0718",	x"071f",	x"06dd",	
												x"0711",	x"0713",	x"0718",	x"06fa",	
												x"0718",	x"0719",	x"0727",	x"0734",	
												x"0726",	x"0723",	x"071a",	x"0718",	
												x"071c",	x"0708",	x"074c",	x"06ea",	
												x"072f",	x"0721",	x"072d",	x"0704",	
												x"0714",	x"0701",	x"0722",	x"0701",	
												x"0751",	x"0710",	x"0746",	x"0720",	
												x"06f7",	x"0720",	x"0004",	x"000a",	
												x"2591",	x"ce46",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"3140",	
												x"06f7",	x"06c8",	x"0705",	x"06f6",	
												x"0707",	x"06f9",	x"070d",	x"0706",	
												x"06e7",	x"06c9",	x"0704",	x"06f1",	
												x"06d6",	x"06af",	x"06d5",	x"06eb",	
												x"071f",	x"06cc",	x"072e",	x"0709",	
												x"072d",	x"06f7",	x"073b",	x"0732",	
												x"073f",	x"06ec",	x"0755",	x"0720",	
												x"0758",	x"0742",	x"073f",	x"0732",	
												x"0766",	x"0737",	x"0770",	x"0752",	
												x"0756",	x"0765",	x"0766",	x"0751",	
												x"076f",	x"0757",	x"0752",	x"073a",	
												x"0770",	x"0742",	x"073e",	x"075d",	
												x"076e",	x"0746",	x"077f",	x"0744",	
												x"0771",	x"075a",	x"0780",	x"0776",	
												x"077c",	x"075d",	x"0798",	x"0769",	
												x"0799",	x"0762",	x"0722",	x"076e",	
												x"5031",	x"3140",	x"0730",	x"072e",	
												x"074b",	x"074c",	x"076b",	x"072e",	
												x"0741",	x"075b",	x"077a",	x"070a",	
												x"074b",	x"072e",	x"071e",	x"0714",	
												x"0727",	x"0720",	x"076c",	x"0722",	
												x"077e",	x"0749",	x"077b",	x"074e",	
												x"0779",	x"073f",	x"0785",	x"0739",	
												x"0787",	x"0751",	x"077e",	x"0767",	
												x"0763",	x"0759",	x"078d",	x"0752",	
												x"0793",	x"0771",	x"0788",	x"0762",	
												x"07a0",	x"075f",	x"07a6",	x"075e",	
												x"07ae",	x"0768",	x"07bc",	x"0769",	
												x"0793",	x"0768",	x"07c0",	x"076b",	
												x"07b8",	x"0779",	x"07d6",	x"0763",	
												x"07b5",	x"077e",	x"07c1",	x"077f",	
												x"07e0",	x"077d",	x"07ca",	x"078c",	
												x"0732",	x"0779",	x"6031",	x"3140",	
												x"074a",	x"0723",	x"0756",	x"0731",	
												x"0762",	x"072f",	x"0747",	x"072d",	
												x"0751",	x"072f",	x"0759",	x"0746",	
												x"0774",	x"070e",	x"074b",	x"0729",	
												x"0778",	x"0705",	x"076b",	x"0739",	
												x"079d",	x"074a",	x"07a2",	x"0775",	
												x"079f",	x"0762",	x"079a",	x"0778",	
												x"07b8",	x"077f",	x"0787",	x"077b",	
												x"07ac",	x"0771",	x"07bb",	x"078f",	
												x"07be",	x"078f",	x"07d6",	x"07b7",	
												x"07c9",	x"0794",	x"07ee",	x"0792",	
												x"07f3",	x"079d",	x"07c0",	x"07b7",	
												x"07e9",	x"0798",	x"07f4",	x"07b3",	
												x"07ce",	x"07b5",	x"080a",	x"079f",	
												x"080a",	x"079d",	x"081b",	x"0797",	
												x"081b",	x"07b0",	x"074e",	x"07ad",	
												x"7031",	x"3140",	x"07a6",	x"0751",	
												x"0784",	x"0770",	x"07c0",	x"0766",	
												x"079a",	x"0768",	x"07a2",	x"0765",	
												x"078e",	x"0762",	x"077f",	x"0781",	
												x"0776",	x"075d",	x"07c4",	x"0757",	
												x"0800",	x"0781",	x"083b",	x"07af",	
												x"0816",	x"07c4",	x"0800",	x"07cc",	
												x"0834",	x"07e9",	x"080a",	x"07e2",	
												x"0828",	x"07f2",	x"0832",	x"07f7",	
												x"0811",	x"07fe",	x"0841",	x"0805",	
												x"084b",	x"0815",	x"0840",	x"0822",	
												x"086f",	x"0825",	x"0861",	x"083a",	
												x"082d",	x"0829",	x"0865",	x"0817",	
												x"0865",	x"0823",	x"0856",	x"082b",	
												x"085c",	x"0839",	x"0868",	x"082d",	
												x"087e",	x"0865",	x"0854",	x"0840",	
												x"0680",	x"085a",	x"0004",	x"000a",	
												x"6db5",	x"0218",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"0241",	
												x"0750",	x"0740",	x"0746",	x"0749",	
												x"0726",	x"073a",	x"075a",	x"072f",	
												x"073d",	x"0754",	x"0749",	x"0748",	
												x"0758",	x"0775",	x"0767",	x"0770",	
												x"079a",	x"078f",	x"07af",	x"07cc",	
												x"0768",	x"0789",	x"0776",	x"0772",	
												x"0780",	x"076e",	x"0784",	x"079b",	
												x"0775",	x"078f",	x"072c",	x"0797",	
												x"0798",	x"0784",	x"078b",	x"079b",	
												x"078d",	x"0779",	x"0787",	x"07a5",	
												x"0750",	x"075f",	x"077e",	x"0760",	
												x"0769",	x"0785",	x"077a",	x"075e",	
												x"0776",	x"07ac",	x"077e",	x"07a6",	
												x"0777",	x"0778",	x"0790",	x"07b3",	
												x"0793",	x"078c",	x"0792",	x"0771",	
												x"07a2",	x"077e",	x"0725",	x"0795",	
												x"102e",	x"0241",	x"0726",	x"073c",	
												x"075d",	x"073e",	x"0706",	x"075d",	
												x"06fe",	x"071e",	x"073b",	x"0745",	
												x"075b",	x"0743",	x"075d",	x"075c",	
												x"0765",	x"076e",	x"0772",	x"0761",	
												x"0796",	x"078a",	x"0759",	x"078a",	
												x"075d",	x"0772",	x"0762",	x"0754",	
												x"077d",	x"078e",	x"077c",	x"0779",	
												x"0757",	x"0777",	x"0767",	x"0756",	
												x"0761",	x"0775",	x"0778",	x"0751",	
												x"0771",	x"0782",	x"077f",	x"076e",	
												x"0774",	x"07aa",	x"0755",	x"078c",	
												x"076c",	x"0759",	x"075b",	x"078b",	
												x"0787",	x"0782",	x"076d",	x"0795",	
												x"0775",	x"0780",	x"077d",	x"077b",	
												x"0765",	x"0775",	x"0783",	x"0784",	
												x"071f",	x"0791",	x"202e",	x"0241",	
												x"072e",	x"0725",	x"0701",	x"072e",	
												x"06f5",	x"0709",	x"0716",	x"072c",	
												x"073c",	x"0766",	x"072e",	x"0732",	
												x"072a",	x"0743",	x"073e",	x"0759",	
												x"076c",	x"0752",	x"075b",	x"076d",	
												x"0742",	x"0759",	x"0751",	x"077c",	
												x"074f",	x"0764",	x"0748",	x"0756",	
												x"073f",	x"0764",	x"0745",	x"0761",	
												x"0754",	x"075b",	x"075d",	x"0763",	
												x"075f",	x"0765",	x"075e",	x"0766",	
												x"0747",	x"073d",	x"0745",	x"0732",	
												x"0755",	x"0746",	x"0743",	x"074a",	
												x"0773",	x"0775",	x"0753",	x"0764",	
												x"0733",	x"075a",	x"076f",	x"0751",	
												x"076d",	x"075d",	x"076d",	x"0758",	
												x"076c",	x"0757",	x"0704",	x"0750",	
												x"302e",	x"0241",	x"0706",	x"06c4",	
												x"071c",	x"070e",	x"06f6",	x"0721",	
												x"0717",	x"06f4",	x"0725",	x"070c",	
												x"0748",	x"0726",	x"0738",	x"0739",	
												x"0712",	x"0735",	x"074b",	x"0718",	
												x"074d",	x"073e",	x"0744",	x"073a",	
												x"0734",	x"075c",	x"0745",	x"0734",	
												x"073f",	x"0761",	x"075a",	x"0761",	
												x"072b",	x"074b",	x"0747",	x"072c",	
												x"074b",	x"073c",	x"0739",	x"074e",	
												x"075a",	x"073c",	x"073c",	x"0746",	
												x"074a",	x"0728",	x"0744",	x"073c",	
												x"073a",	x"074d",	x"077c",	x"074b",	
												x"0777",	x"0752",	x"075f",	x"072e",	
												x"077c",	x"075c",	x"075c",	x"0758",	
												x"0765",	x"0742",	x"0781",	x"0760",	
												x"0704",	x"0764",	x"0004",	x"000a",	
												x"4a87",	x"3b72",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"0242",	
												x"072d",	x"070b",	x"073a",	x"0708",	
												x"0726",	x"0715",	x"072b",	x"070a",	
												x"071a",	x"071f",	x"072d",	x"0734",	
												x"0735",	x"0739",	x"0724",	x"0744",	
												x"0765",	x"073f",	x"0761",	x"0773",	
												x"074f",	x"075a",	x"0759",	x"0752",	
												x"0765",	x"074c",	x"075f",	x"075e",	
												x"0771",	x"0752",	x"0759",	x"076c",	
												x"0771",	x"0761",	x"0784",	x"0777",	
												x"0785",	x"0778",	x"0782",	x"0778",	
												x"078b",	x"0794",	x"0790",	x"077f",	
												x"0789",	x"0784",	x"0764",	x"0796",	
												x"07aa",	x"07a0",	x"0787",	x"0773",	
												x"078d",	x"077f",	x"079d",	x"0796",	
												x"07a8",	x"0783",	x"07aa",	x"0780",	
												x"07ad",	x"0791",	x"0750",	x"077e",	
												x"502e",	x"0242",	x"0768",	x"0736",	
												x"078a",	x"0748",	x"0765",	x"075c",	
												x"076f",	x"0751",	x"076f",	x"074f",	
												x"07a0",	x"0787",	x"07b1",	x"078c",	
												x"0782",	x"078b",	x"0797",	x"078a",	
												x"0792",	x"0784",	x"07a3",	x"0796",	
												x"07a6",	x"07a8",	x"07aa",	x"07a7",	
												x"0781",	x"079b",	x"07c0",	x"0794",	
												x"07a7",	x"0799",	x"07c1",	x"0798",	
												x"07b1",	x"07b6",	x"07a7",	x"0780",	
												x"07a1",	x"079d",	x"07c8",	x"078e",	
												x"07bd",	x"07a6",	x"07c7",	x"0789",	
												x"07c0",	x"07b1",	x"07d3",	x"07b6",	
												x"07c6",	x"0797",	x"07cf",	x"079b",	
												x"07da",	x"0788",	x"07ca",	x"07a3",	
												x"07f7",	x"07aa",	x"07f3",	x"07b7",	
												x"076b",	x"07b4",	x"602e",	x"0242",	
												x"0784",	x"0730",	x"075c",	x"0759",	
												x"0780",	x"075a",	x"078e",	x"075a",	
												x"0771",	x"0767",	x"078b",	x"074b",	
												x"07a8",	x"0773",	x"07b0",	x"0787",	
												x"07c1",	x"078e",	x"07be",	x"07ba",	
												x"07e1",	x"07ae",	x"07e2",	x"07b1",	
												x"07cf",	x"07ab",	x"0805",	x"07ba",	
												x"07f3",	x"07bd",	x"07cd",	x"07db",	
												x"07eb",	x"07cb",	x"07ee",	x"07df",	
												x"07e2",	x"07d3",	x"07fd",	x"07c5",	
												x"07ff",	x"07c8",	x"07f4",	x"07e7",	
												x"07e6",	x"07f0",	x"07f2",	x"07f5",	
												x"081c",	x"07d2",	x"07f2",	x"07e8",	
												x"0804",	x"07ce",	x"082e",	x"07dc",	
												x"0825",	x"07d4",	x"0829",	x"0806",	
												x"0829",	x"07e4",	x"079c",	x"07f2",	
												x"702e",	x"0242",	x"07c3",	x"0783",	
												x"07b5",	x"07a0",	x"07dd",	x"07a0",	
												x"07dc",	x"07c6",	x"07bd",	x"07cc",	
												x"07f4",	x"07ce",	x"07fb",	x"0818",	
												x"07ee",	x"07ee",	x"081e",	x"07e2",	
												x"0831",	x"07f4",	x"082e",	x"0813",	
												x"0841",	x"081e",	x"0843",	x"0818",	
												x"0835",	x"0833",	x"082d",	x"082d",	
												x"0836",	x"0844",	x"085e",	x"0818",	
												x"0874",	x"0841",	x"087d",	x"084e",	
												x"0885",	x"0852",	x"084f",	x"0843",	
												x"0880",	x"0846",	x"0864",	x"085f",	
												x"0836",	x"0857",	x"086c",	x"0859",	
												x"08b7",	x"0881",	x"0889",	x"086d",	
												x"08c7",	x"0862",	x"08bd",	x"0887",	
												x"08cd",	x"088f",	x"08ac",	x"0893",	
												x"05d3",	x"089d",	x"0004",	x"000a",	
												x"82d4",	x"664d",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"1243",	
												x"05d8",	x"05e0",	x"05f5",	x"05d7",	
												x"05ea",	x"05fe",	x"05e8",	x"05fe",	
												x"05e3",	x"05f4",	x"0611",	x"05e2",	
												x"05df",	x"0621",	x"05cf",	x"05ec",	
												x"0611",	x"0605",	x"061f",	x"0609",	
												x"0628",	x"0614",	x"062d",	x"061e",	
												x"060c",	x"0653",	x"0634",	x"0616",	
												x"05ee",	x"0639",	x"05d8",	x"0610",	
												x"061c",	x"0605",	x"0612",	x"063e",	
												x"0621",	x"0610",	x"0629",	x"063c",	
												x"060a",	x"0628",	x"0617",	x"061d",	
												x"0613",	x"0609",	x"0605",	x"0618",	
												x"0620",	x"0606",	x"0632",	x"0613",	
												x"062e",	x"0628",	x"0620",	x"0614",	
												x"061b",	x"0618",	x"0621",	x"0624",	
												x"0636",	x"0601",	x"05e1",	x"060b",	
												x"102e",	x"1243",	x"05cc",	x"05ce",	
												x"05c8",	x"05d0",	x"05df",	x"05cc",	
												x"05e8",	x"05e8",	x"05e4",	x"05e7",	
												x"05f8",	x"05e7",	x"05ee",	x"05e7",	
												x"05d0",	x"0601",	x"0606",	x"05ef",	
												x"0614",	x"060e",	x"060f",	x"0611",	
												x"0606",	x"061a",	x"0610",	x"061f",	
												x"0619",	x"0611",	x"05f7",	x"0627",	
												x"05b8",	x"05fb",	x"05f7",	x"05fb",	
												x"05fb",	x"0628",	x"05f9",	x"0612",	
												x"0609",	x"0607",	x"05fc",	x"0615",	
												x"05fb",	x"0610",	x"060c",	x"060c",	
												x"05f0",	x"0618",	x"061a",	x"05fd",	
												x"0617",	x"060d",	x"061a",	x"0613",	
												x"0632",	x"0616",	x"062a",	x"061f",	
												x"0627",	x"0630",	x"061b",	x"0623",	
												x"05b8",	x"061b",	x"202e",	x"1243",	
												x"05b2",	x"05b1",	x"05cf",	x"05d1",	
												x"05ca",	x"05d5",	x"05ce",	x"05df",	
												x"05eb",	x"05e4",	x"05e5",	x"05fb",	
												x"05e8",	x"05f9",	x"05d9",	x"05fc",	
												x"05dd",	x"0608",	x"05e9",	x"05fe",	
												x"0600",	x"0605",	x"05f4",	x"05f3",	
												x"05fc",	x"05f1",	x"05f8",	x"05fd",	
												x"05f4",	x"0605",	x"05ce",	x"05f7",	
												x"05f1",	x"05e2",	x"05e6",	x"05fc",	
												x"0604",	x"0601",	x"05f7",	x"061d",	
												x"05ff",	x"05e5",	x"05fc",	x"05fb",	
												x"05f8",	x"05f6",	x"05dc",	x"05fc",	
												x"05e3",	x"05df",	x"0616",	x"0601",	
												x"0606",	x"0600",	x"060d",	x"05fb",	
												x"0617",	x"0600",	x"060d",	x"0615",	
												x"060d",	x"05fa",	x"05c7",	x"05f0",	
												x"302e",	x"1243",	x"05c7",	x"05a6",	
												x"059d",	x"059d",	x"05b2",	x"05aa",	
												x"05c9",	x"05bd",	x"05c5",	x"05e0",	
												x"05c6",	x"05c4",	x"05e0",	x"05c0",	
												x"05a9",	x"05ca",	x"05e7",	x"05da",	
												x"05e3",	x"05db",	x"05fa",	x"05d4",	
												x"05f8",	x"05ee",	x"05f0",	x"05f2",	
												x"05f0",	x"05eb",	x"05f4",	x"05e6",	
												x"05c0",	x"05dd",	x"05fd",	x"05d8",	
												x"05ee",	x"05f4",	x"060f",	x"05f0",	
												x"0606",	x"05fd",	x"05fc",	x"0604",	
												x"060a",	x"05fe",	x"05f5",	x"05f4",	
												x"05f4",	x"05eb",	x"0605",	x"05f7",	
												x"060f",	x"05f4",	x"0615",	x"0611",	
												x"0617",	x"060b",	x"0618",	x"05fb",	
												x"0616",	x"0600",	x"061f",	x"05fd",	
												x"05d0",	x"0604",	x"0004",	x"000a",	
												x"9bd6",	x"cb01",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"1244",	
												x"05e0",	x"05b0",	x"05db",	x"05c9",	
												x"05e1",	x"05c5",	x"0602",	x"05e2",	
												x"05c1",	x"05d4",	x"05da",	x"05e4",	
												x"05da",	x"05de",	x"05f1",	x"05eb",	
												x"05f0",	x"05ee",	x"0607",	x"061c",	
												x"060f",	x"0619",	x"0609",	x"0615",	
												x"060a",	x"05f9",	x"05fe",	x"0603",	
												x"0605",	x"05f7",	x"0613",	x"0607",	
												x"0617",	x"05da",	x"061e",	x"0610",	
												x"0627",	x"062a",	x"061c",	x"062a",	
												x"062f",	x"0630",	x"061a",	x"062a",	
												x"0625",	x"0616",	x"0604",	x"0628",	
												x"0634",	x"0632",	x"063e",	x"0631",	
												x"0635",	x"061f",	x"0655",	x"0647",	
												x"063e",	x"0645",	x"065e",	x"0642",	
												x"0652",	x"0663",	x"05ff",	x"0635",	
												x"502e",	x"1244",	x"0612",	x"05e7",	
												x"0602",	x"05f7",	x"0623",	x"05f4",	
												x"0626",	x"061a",	x"0624",	x"0622",	
												x"0620",	x"05f2",	x"0648",	x"0609",	
												x"061a",	x"063a",	x"063f",	x"05fe",	
												x"0642",	x"062f",	x"0646",	x"062d",	
												x"065f",	x"0641",	x"0650",	x"0642",	
												x"063d",	x"063f",	x"063c",	x"063c",	
												x"062b",	x"062a",	x"0650",	x"0617",	
												x"064a",	x"0652",	x"0650",	x"0637",	
												x"0666",	x"0643",	x"0659",	x"0640",	
												x"0668",	x"0642",	x"066d",	x"0625",	
												x"0657",	x"064a",	x"0644",	x"0649",	
												x"0682",	x"064e",	x"0675",	x"064f",	
												x"0688",	x"065c",	x"067a",	x"0651",	
												x"0687",	x"0662",	x"068b",	x"0663",	
												x"0635",	x"0652",	x"602e",	x"1244",	
												x"0612",	x"05eb",	x"0611",	x"05ee",	
												x"0626",	x"05ed",	x"062d",	x"061a",	
												x"0640",	x"0621",	x"063d",	x"0603",	
												x"0649",	x"063a",	x"0638",	x"0626",	
												x"0659",	x"0617",	x"0673",	x"0646",	
												x"0664",	x"064b",	x"0667",	x"0654",	
												x"0679",	x"0651",	x"0665",	x"0668",	
												x"0661",	x"064b",	x"0658",	x"0658",	
												x"066a",	x"065a",	x"067a",	x"0670",	
												x"0685",	x"0662",	x"06a4",	x"0669",	
												x"0697",	x"0697",	x"0692",	x"0677",	
												x"0698",	x"066d",	x"0674",	x"0680",	
												x"069d",	x"0678",	x"069e",	x"067c",	
												x"06b4",	x"068c",	x"06b2",	x"0685",	
												x"0693",	x"0676",	x"06a6",	x"067a",	
												x"06bd",	x"068a",	x"0650",	x"0669",	
												x"702e",	x"1244",	x"0652",	x"0616",	
												x"0640",	x"0632",	x"0644",	x"0624",	
												x"0687",	x"0626",	x"068e",	x"062e",	
												x"0679",	x"065e",	x"0671",	x"0665",	
												x"068e",	x"0664",	x"06a5",	x"065d",	
												x"06ca",	x"0696",	x"06ae",	x"06a8",	
												x"06bd",	x"069f",	x"06b7",	x"06bb",	
												x"06dd",	x"06bb",	x"06b4",	x"069a",	
												x"0698",	x"06a1",	x"06cc",	x"06ad",	
												x"06db",	x"06c9",	x"06d3",	x"06b5",	
												x"06e0",	x"06b3",	x"06f3",	x"06d4",	
												x"06ed",	x"06ef",	x"06dc",	x"06c5",	
												x"06d0",	x"06c3",	x"06e3",	x"06dc",	
												x"06fc",	x"06cf",	x"06f3",	x"06f1",	
												x"072d",	x"06fd",	x"0732",	x"06fc",	
												x"071e",	x"0702",	x"070a",	x"0706",	
												x"06d6",	x"06ed",	x"0004",	x"000a",	
												x"d10d",	x"f38c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"2245",	
												x"06ba",	x"06cd",	x"06d2",	x"06b3",	
												x"06e9",	x"06f0",	x"06ee",	x"06fa",	
												x"06eb",	x"06e1",	x"06e6",	x"06ed",	
												x"070a",	x"06fe",	x"06fc",	x"06fa",	
												x"06ee",	x"06f8",	x"0709",	x"072f",	
												x"06f2",	x"0725",	x"0723",	x"0729",	
												x"06f7",	x"0704",	x"0707",	x"0738",	
												x"06fd",	x"0719",	x"06d5",	x"0708",	
												x"06e6",	x"06df",	x"06f3",	x"06fb",	
												x"06d7",	x"06ee",	x"070e",	x"0704",	
												x"071e",	x"0742",	x"06d6",	x"0725",	
												x"06d9",	x"06e0",	x"06e9",	x"06e7",	
												x"06de",	x"06f2",	x"0709",	x"06f5",	
												x"06e7",	x"06e8",	x"06f6",	x"06f8",	
												x"072b",	x"06ee",	x"073f",	x"0717",	
												x"070e",	x"0707",	x"06a8",	x"06f8",	
												x"102e",	x"2245",	x"0690",	x"0691",	
												x"06c6",	x"06a8",	x"06a5",	x"06d2",	
												x"06ad",	x"06bf",	x"06cf",	x"06da",	
												x"06d0",	x"06d0",	x"06d1",	x"06e1",	
												x"06de",	x"06b5",	x"06eb",	x"06c9",	
												x"06f6",	x"06fb",	x"06fe",	x"06fd",	
												x"06f0",	x"06fb",	x"06ed",	x"06fc",	
												x"06e7",	x"06eb",	x"06e0",	x"06f1",	
												x"0691",	x"06ee",	x"06d6",	x"06c1",	
												x"06e9",	x"06e3",	x"06fa",	x"06fc",	
												x"06fc",	x"070a",	x"06f3",	x"0702",	
												x"06e6",	x"06fb",	x"06e6",	x"06f2",	
												x"06b6",	x"06ee",	x"06ec",	x"0706",	
												x"06f6",	x"06fb",	x"06f9",	x"06fa",	
												x"0719",	x"071a",	x"0710",	x"070b",	
												x"070b",	x"0711",	x"0707",	x"0709",	
												x"068e",	x"0702",	x"202e",	x"2245",	
												x"0694",	x"068a",	x"06a4",	x"069f",	
												x"069d",	x"069e",	x"069c",	x"06b8",	
												x"06b7",	x"06cb",	x"06a7",	x"06be",	
												x"06b7",	x"06ca",	x"06b1",	x"06d3",	
												x"06e5",	x"06d4",	x"06d6",	x"06fd",	
												x"06d6",	x"06fb",	x"06d4",	x"06e8",	
												x"06c0",	x"06ea",	x"06d5",	x"06e3",	
												x"06d3",	x"06df",	x"06ad",	x"06d7",	
												x"06b8",	x"06c1",	x"06c3",	x"06b6",	
												x"06df",	x"06c9",	x"06ce",	x"06d9",	
												x"06ea",	x"06d6",	x"06e5",	x"06fb",	
												x"06da",	x"06e7",	x"06bc",	x"06cf",	
												x"06c6",	x"06cf",	x"06e4",	x"06ea",	
												x"06d1",	x"06ea",	x"06f6",	x"06dd",	
												x"06d3",	x"06c8",	x"06ed",	x"06d9",	
												x"06e8",	x"06ed",	x"0667",	x"06d5",	
												x"302e",	x"2245",	x"0678",	x"0658",	
												x"068c",	x"0676",	x"0699",	x"0687",	
												x"06a1",	x"068f",	x"06ae",	x"0696",	
												x"069c",	x"06a4",	x"06ac",	x"06c3",	
												x"0691",	x"06bc",	x"06af",	x"06ab",	
												x"06c3",	x"06b8",	x"06ca",	x"06d3",	
												x"06cf",	x"06c8",	x"06c2",	x"06cf",	
												x"06ca",	x"06c2",	x"06c2",	x"06bc",	
												x"0691",	x"06b5",	x"06a7",	x"068b",	
												x"06b9",	x"069f",	x"06ab",	x"06a5",	
												x"06bf",	x"06c5",	x"06d1",	x"06b8",	
												x"06d2",	x"06dd",	x"06da",	x"06d5",	
												x"06c9",	x"06d9",	x"06e5",	x"06d0",	
												x"06cf",	x"06c9",	x"06eb",	x"06d6",	
												x"06ed",	x"06d1",	x"06f6",	x"06cd",	
												x"06f5",	x"06c8",	x"06f0",	x"06d2",	
												x"0672",	x"06cc",	x"0004",	x"000a",	
												x"0a30",	x"7b5f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"2246",	
												x"0693",	x"0689",	x"06aa",	x"069c",	
												x"06a1",	x"06ca",	x"06ac",	x"06cb",	
												x"06bc",	x"06ae",	x"06c0",	x"06b6",	
												x"06ce",	x"06db",	x"06b7",	x"06b7",	
												x"06dd",	x"06c7",	x"06e0",	x"06e9",	
												x"06cc",	x"06e9",	x"06d0",	x"06e1",	
												x"06da",	x"06dc",	x"06ec",	x"06e7",	
												x"06fa",	x"0710",	x"06d5",	x"0705",	
												x"06fb",	x"06ea",	x"06f5",	x"0700",	
												x"06f7",	x"06f6",	x"0703",	x"06f2",	
												x"0703",	x"06ed",	x"072e",	x"070a",	
												x"0722",	x"0713",	x"06e8",	x"06fc",	
												x"071b",	x"0705",	x"0727",	x"070c",	
												x"0727",	x"0721",	x"0731",	x"0715",	
												x"072b",	x"071a",	x"0727",	x"0713",	
												x"073f",	x"0710",	x"06ae",	x"070f",	
												x"502e",	x"2246",	x"06f4",	x"069f",	
												x"06da",	x"06d2",	x"06ad",	x"06e7",	
												x"06ce",	x"06b7",	x"06f9",	x"06e9",	
												x"06ec",	x"06f8",	x"06fe",	x"06f1",	
												x"06f1",	x"0704",	x"071c",	x"06f8",	
												x"0732",	x"071f",	x"0721",	x"0700",	
												x"0716",	x"0728",	x"0713",	x"071c",	
												x"070f",	x"0715",	x"0723",	x"0701",	
												x"06e0",	x"070c",	x"06f9",	x"06f2",	
												x"071b",	x"070e",	x"0721",	x"0711",	
												x"0728",	x"0714",	x"0725",	x"070f",	
												x"0741",	x"0726",	x"071e",	x"071e",	
												x"0733",	x"071d",	x"074d",	x"0726",	
												x"074e",	x"0735",	x"0758",	x"0719",	
												x"075a",	x"0720",	x"076a",	x"0730",	
												x"076a",	x"073f",	x"075f",	x"0732",	
												x"06c3",	x"0734",	x"602e",	x"2246",	
												x"06f8",	x"06a5",	x"06e8",	x"06b5",	
												x"06ed",	x"06e9",	x"070d",	x"06f0",	
												x"071d",	x"06ea",	x"0722",	x"070c",	
												x"0728",	x"0711",	x"071b",	x"0722",	
												x"0755",	x"0712",	x"0723",	x"0751",	
												x"0720",	x"072a",	x"0759",	x"0725",	
												x"0753",	x"073c",	x"0769",	x"0744",	
												x"0750",	x"0731",	x"071f",	x"0743",	
												x"073a",	x"071f",	x"0747",	x"0752",	
												x"0766",	x"0746",	x"0764",	x"0753",	
												x"0763",	x"076d",	x"0771",	x"0762",	
												x"0767",	x"0764",	x"076f",	x"0765",	
												x"0775",	x"0745",	x"0793",	x"074c",	
												x"07a6",	x"0755",	x"07af",	x"0779",	
												x"0797",	x"0784",	x"07a5",	x"076f",	
												x"07a4",	x"077a",	x"0719",	x"0779",	
												x"702e",	x"2246",	x"0724",	x"070c",	
												x"0712",	x"070a",	x"071b",	x"0715",	
												x"0755",	x"0712",	x"0724",	x"071f",	
												x"0766",	x"0734",	x"0748",	x"0762",	
												x"0755",	x"0744",	x"0783",	x"076d",	
												x"078f",	x"0790",	x"0785",	x"0784",	
												x"0790",	x"07a7",	x"0786",	x"0797",	
												x"07cc",	x"0786",	x"0795",	x"07a3",	
												x"0794",	x"07b8",	x"07bd",	x"0785",	
												x"07cf",	x"07b4",	x"07eb",	x"078d",	
												x"0808",	x"0807",	x"07c6",	x"07bd",	
												x"07ce",	x"07c8",	x"07d4",	x"07b1",	
												x"07d9",	x"07c1",	x"07c6",	x"07de",	
												x"07f1",	x"07c9",	x"07ec",	x"07cf",	
												x"07cd",	x"07d8",	x"0821",	x"07da",	
												x"082b",	x"080b",	x"0811",	x"0804",	
												x"06d9",	x"080b",	x"0004",	x"000a",	
												x"3dc1",	x"a59a",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"3247",	
												x"06d4",	x"06d6",	x"06fe",	x"06fc",	
												x"06ac",	x"06c8",	x"06bc",	x"06c2",	
												x"06f0",	x"06d6",	x"070e",	x"0706",	
												x"0703",	x"0722",	x"06e6",	x"0700",	
												x"0722",	x"0717",	x"0725",	x"0737",	
												x"06f1",	x"0718",	x"0719",	x"0736",	
												x"0703",	x"0723",	x"072b",	x"071b",	
												x"06fa",	x"0719",	x"06e2",	x"070e",	
												x"06fa",	x"0700",	x"0704",	x"0722",	
												x"0712",	x"070f",	x"0702",	x"0712",	
												x"0711",	x"06fe",	x"073b",	x"0724",	
												x"072e",	x"0734",	x"06f5",	x"0739",	
												x"0701",	x"06ef",	x"0707",	x"070a",	
												x"0708",	x"0706",	x"0725",	x"0717",	
												x"070e",	x"0714",	x"0728",	x"0718",	
												x"0706",	x"072a",	x"06dc",	x"071e",	
												x"102e",	x"3247",	x"06af",	x"06bf",	
												x"06c4",	x"06b8",	x"06c8",	x"06bc",	
												x"06d4",	x"06e2",	x"06da",	x"06d1",	
												x"06f1",	x"06d8",	x"06e0",	x"06f2",	
												x"06f2",	x"06ea",	x"06ff",	x"06fc",	
												x"0713",	x"070a",	x"06ed",	x"071f",	
												x"070b",	x"06ec",	x"06c9",	x"070e",	
												x"06e3",	x"06dd",	x"06eb",	x"06ea",	
												x"06a6",	x"06f3",	x"06d1",	x"06de",	
												x"06d2",	x"06e4",	x"06f1",	x"06bd",	
												x"0714",	x"0702",	x"06ea",	x"0706",	
												x"06f2",	x"06fb",	x"070f",	x"06ff",	
												x"06d5",	x"0702",	x"06ee",	x"06ea",	
												x"070d",	x"06f8",	x"06db",	x"06ef",	
												x"070e",	x"06ed",	x"070c",	x"070b",	
												x"0726",	x"0729",	x"0735",	x"0736",	
												x"06da",	x"0730",	x"202e",	x"3247",	
												x"06a8",	x"06d0",	x"069f",	x"06c6",	
												x"06af",	x"06ac",	x"06d4",	x"06d9",	
												x"06d0",	x"06de",	x"06d5",	x"070a",	
												x"06de",	x"070a",	x"06bc",	x"06fb",	
												x"06f4",	x"06f6",	x"06f3",	x"0710",	
												x"06e3",	x"070c",	x"06f2",	x"0707",	
												x"06db",	x"06fa",	x"06eb",	x"06f6",	
												x"06d5",	x"06e7",	x"06b1",	x"06dc",	
												x"06da",	x"06c1",	x"06db",	x"06ea",	
												x"06d8",	x"06c4",	x"06e4",	x"06e2",	
												x"06f9",	x"06c2",	x"06f7",	x"06dc",	
												x"06e7",	x"06f2",	x"06d4",	x"06df",	
												x"06e0",	x"06f7",	x"06e2",	x"06e4",	
												x"06e7",	x"06ef",	x"06ff",	x"06f6",	
												x"06f5",	x"06ff",	x"0702",	x"06e4",	
												x"06f0",	x"06ea",	x"0690",	x"06df",	
												x"302e",	x"3247",	x"0684",	x"068d",	
												x"069e",	x"069b",	x"06a0",	x"068a",	
												x"06a9",	x"06c1",	x"06ac",	x"06ba",	
												x"06ba",	x"06b0",	x"06b1",	x"06af",	
												x"06a1",	x"06bd",	x"06cf",	x"06d0",	
												x"06b3",	x"06cb",	x"06dd",	x"06cb",	
												x"06cd",	x"06d9",	x"06c1",	x"06cf",	
												x"06a3",	x"06ad",	x"06bc",	x"06a9",	
												x"0696",	x"06bc",	x"06c5",	x"06bb",	
												x"06b9",	x"06b9",	x"06c0",	x"06ba",	
												x"06e6",	x"06d7",	x"06ec",	x"06c6",	
												x"06d7",	x"06db",	x"06e6",	x"06d5",	
												x"06ba",	x"06e3",	x"06de",	x"06c9",	
												x"06ea",	x"06d9",	x"06e0",	x"06de",	
												x"06f4",	x"06d3",	x"06fc",	x"06e0",	
												x"0700",	x"06df",	x"06ee",	x"06e7",	
												x"06b4",	x"06cd",	x"0004",	x"000a",	
												x"1170",	x"c29d",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"3248",	
												x"067e",	x"0685",	x"06dc",	x"0690",	
												x"06a3",	x"06ae",	x"06b3",	x"06b3",	
												x"06b6",	x"06c0",	x"06c2",	x"06ba",	
												x"06bc",	x"06e4",	x"06b1",	x"06f5",	
												x"06d4",	x"06e6",	x"06f5",	x"06e5",	
												x"06f6",	x"0709",	x"06e7",	x"0707",	
												x"06fa",	x"06d3",	x"06fb",	x"06f6",	
												x"06db",	x"06ef",	x"06db",	x"06f4",	
												x"06f9",	x"06de",	x"06f2",	x"06f7",	
												x"0702",	x"0713",	x"070b",	x"0728",	
												x"0708",	x"06f2",	x"0709",	x"0708",	
												x"071a",	x"0710",	x"0707",	x"071a",	
												x"070b",	x"0724",	x"0706",	x"0709",	
												x"071b",	x"0712",	x"072d",	x"0725",	
												x"072c",	x"071e",	x"0731",	x"0714",	
												x"0722",	x"0717",	x"06db",	x"0728",	
												x"502e",	x"3248",	x"06d0",	x"06ba",	
												x"06da",	x"06e2",	x"06c9",	x"06b9",	
												x"06e5",	x"06c3",	x"06fc",	x"06d2",	
												x"0703",	x"0717",	x"0723",	x"072b",	
												x"0705",	x"0729",	x"0719",	x"071b",	
												x"0727",	x"0711",	x"073c",	x"0719",	
												x"072a",	x"0737",	x"073a",	x"071a",	
												x"070c",	x"071f",	x"0704",	x"0701",	
												x"0701",	x"0719",	x"072a",	x"0717",	
												x"071e",	x"0737",	x"073c",	x"070d",	
												x"0738",	x"0727",	x"0748",	x"0715",	
												x"0753",	x"072f",	x"0760",	x"073a",	
												x"0721",	x"0734",	x"0740",	x"0722",	
												x"0750",	x"0721",	x"0753",	x"0725",	
												x"0775",	x"0735",	x"0777",	x"0758",	
												x"0761",	x"0738",	x"0756",	x"0738",	
												x"06cd",	x"0716",	x"602e",	x"3248",	
												x"06e4",	x"06b4",	x"06dc",	x"06f9",	
												x"06f2",	x"06ac",	x"06f6",	x"06d0",	
												x"06f6",	x"06d1",	x"071e",	x"0708",	
												x"072e",	x"072c",	x"0726",	x"071e",	
												x"0737",	x"070b",	x"0753",	x"0739",	
												x"074b",	x"0739",	x"073b",	x"0740",	
												x"072d",	x"0723",	x"072d",	x"0725",	
												x"0740",	x"072b",	x"0734",	x"0735",	
												x"075e",	x"0738",	x"0762",	x"0764",	
												x"0757",	x"074a",	x"076a",	x"073a",	
												x"075f",	x"074e",	x"077a",	x"075d",	
												x"0789",	x"0752",	x"074b",	x"0767",	
												x"0761",	x"0761",	x"0776",	x"0760",	
												x"0783",	x"0758",	x"07ab",	x"077e",	
												x"07b8",	x"0780",	x"0797",	x"0785",	
												x"079b",	x"076e",	x"0722",	x"0772",	
												x"702e",	x"3248",	x"06f7",	x"0725",	
												x"06fc",	x"06fc",	x"0735",	x"06f7",	
												x"0764",	x"072e",	x"074e",	x"074e",	
												x"0757",	x"073d",	x"0748",	x"0760",	
												x"0765",	x"074e",	x"0786",	x"0759",	
												x"07da",	x"07b1",	x"0792",	x"0795",	
												x"07af",	x"0782",	x"07a0",	x"0790",	
												x"07c2",	x"0795",	x"07a9",	x"07a8",	
												x"077b",	x"07b9",	x"0791",	x"0791",	
												x"07b9",	x"079b",	x"07b9",	x"07a7",	
												x"07e7",	x"07c3",	x"07e7",	x"07de",	
												x"07e3",	x"07dc",	x"07d7",	x"07dc",	
												x"07cb",	x"07f3",	x"07e0",	x"07d0",	
												x"07e5",	x"07e3",	x"07ea",	x"07fd",	
												x"0827",	x"080f",	x"0834",	x"0813",	
												x"0835",	x"0815",	x"0807",	x"083a",	
												x"07b6",	x"0803",	x"0004",	x"000a",	
												x"4076",	x"e956",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"0249",	
												x"07bf",	x"07a6",	x"07b8",	x"0795",	
												x"0791",	x"07a3",	x"0799",	x"0796",	
												x"078f",	x"0797",	x"07ad",	x"077a",	
												x"0785",	x"07a8",	x"0726",	x"079f",	
												x"0758",	x"0753",	x"0767",	x"075a",	
												x"0736",	x"0778",	x"0748",	x"0754",	
												x"0762",	x"0757",	x"0795",	x"0790",	
												x"076e",	x"079c",	x"0749",	x"07a3",	
												x"078d",	x"0778",	x"0797",	x"079b",	
												x"079a",	x"07a8",	x"07a7",	x"07b4",	
												x"077e",	x"078f",	x"0790",	x"0784",	
												x"0794",	x"0779",	x"0778",	x"077b",	
												x"077e",	x"0792",	x"078e",	x"07a9",	
												x"07a3",	x"078a",	x"0772",	x"07bf",	
												x"077f",	x"0777",	x"077e",	x"0764",	
												x"07a8",	x"076c",	x"0783",	x"077d",	
												x"102f",	x"0249",	x"077e",	x"07ab",	
												x"076d",	x"0790",	x"0791",	x"0782",	
												x"0779",	x"07a8",	x"0757",	x"0794",	
												x"077a",	x"0773",	x"074c",	x"0778",	
												x"071f",	x"073f",	x"0759",	x"0724",	
												x"0758",	x"0752",	x"0719",	x"074f",	
												x"0746",	x"0742",	x"0731",	x"073e",	
												x"0777",	x"073e",	x"074a",	x"0759",	
												x"0762",	x"075a",	x"0770",	x"074e",	
												x"0774",	x"0771",	x"0789",	x"0771",	
												x"0795",	x"0784",	x"075e",	x"07aa",	
												x"07a2",	x"078d",	x"0798",	x"07bd",	
												x"077d",	x"0781",	x"0777",	x"0794",	
												x"077f",	x"0777",	x"0792",	x"076e",	
												x"0796",	x"0781",	x"07a2",	x"07a2",	
												x"0786",	x"078f",	x"077f",	x"077f",	
												x"0757",	x"078a",	x"202f",	x"0249",	
												x"075b",	x"0769",	x"076c",	x"076a",	
												x"076c",	x"0771",	x"0759",	x"0798",	
												x"0762",	x"0749",	x"073f",	x"0765",	
												x"0768",	x"074d",	x"072a",	x"0785",	
												x"0743",	x"0739",	x"0723",	x"075a",	
												x"06fd",	x"0727",	x"0723",	x"0748",	
												x"0745",	x"0739",	x"0741",	x"076c",	
												x"0742",	x"0761",	x"074b",	x"0769",	
												x"0780",	x"0763",	x"0768",	x"076e",	
												x"076e",	x"075f",	x"0763",	x"076a",	
												x"076a",	x"0744",	x"0770",	x"0763",	
												x"077c",	x"076e",	x"072b",	x"0769",	
												x"0761",	x"0757",	x"0769",	x"076e",	
												x"076b",	x"0776",	x"0777",	x"0773",	
												x"075b",	x"0775",	x"0769",	x"074e",	
												x"0773",	x"0773",	x"0748",	x"075f",	
												x"302f",	x"0249",	x"076c",	x"074b",	
												x"075f",	x"077c",	x"0768",	x"075d",	
												x"0758",	x"073d",	x"074f",	x"0742",	
												x"074d",	x"0743",	x"0762",	x"074b",	
												x"072f",	x"0738",	x"072a",	x"070e",	
												x"0722",	x"072c",	x"071e",	x"070b",	
												x"0710",	x"071c",	x"0743",	x"0726",	
												x"0742",	x"074c",	x"0749",	x"0751",	
												x"0740",	x"0748",	x"073c",	x"0748",	
												x"0759",	x"0750",	x"0756",	x"0755",	
												x"075c",	x"0758",	x"0750",	x"0760",	
												x"075d",	x"0742",	x"0766",	x"074b",	
												x"0742",	x"0749",	x"075a",	x"0742",	
												x"076a",	x"0754",	x"075c",	x"0741",	
												x"075f",	x"076f",	x"075d",	x"0748",	
												x"0760",	x"0743",	x"078f",	x"0748",	
												x"0752",	x"075d",	x"0004",	x"000a",	
												x"5251",	x"41e0",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"024a",	
												x"074c",	x"0745",	x"0756",	x"0726",	
												x"0751",	x"073a",	x"0775",	x"074b",	
												x"0750",	x"074d",	x"077a",	x"074c",	
												x"073e",	x"0753",	x"0741",	x"074d",	
												x"0755",	x"073b",	x"0747",	x"0748",	
												x"074d",	x"075c",	x"0766",	x"0752",	
												x"0771",	x"074b",	x"077d",	x"0767",	
												x"076d",	x"076e",	x"0777",	x"0787",	
												x"078b",	x"0771",	x"07b0",	x"0792",	
												x"07a9",	x"078a",	x"0790",	x"07a6",	
												x"0776",	x"07ae",	x"0798",	x"0779",	
												x"0787",	x"07a7",	x"076f",	x"078a",	
												x"07ae",	x"0789",	x"079f",	x"079c",	
												x"079c",	x"07a0",	x"0799",	x"07a8",	
												x"07ab",	x"0786",	x"07b1",	x"078d",	
												x"07b0",	x"078e",	x"07a2",	x"078f",	
												x"502f",	x"024a",	x"07b2",	x"077c",	
												x"07b2",	x"079d",	x"07b9",	x"07b6",	
												x"07b9",	x"07b0",	x"079f",	x"0786",	
												x"079b",	x"077f",	x"079b",	x"078d",	
												x"0793",	x"0790",	x"0789",	x"078f",	
												x"0792",	x"0780",	x"0763",	x"0788",	
												x"07ac",	x"076f",	x"07af",	x"0794",	
												x"07b1",	x"0797",	x"07ab",	x"07a2",	
												x"07b7",	x"0798",	x"07c4",	x"0794",	
												x"07b1",	x"07ad",	x"07a9",	x"0779",	
												x"07c2",	x"0799",	x"07d8",	x"07bb",	
												x"07df",	x"07b5",	x"07e0",	x"07b1",	
												x"07cc",	x"07b3",	x"07d4",	x"07a3",	
												x"07ea",	x"07aa",	x"07c9",	x"07ba",	
												x"07ce",	x"079c",	x"07d9",	x"078f",	
												x"07ef",	x"079f",	x"07eb",	x"07bf",	
												x"07bf",	x"07bb",	x"602f",	x"024a",	
												x"07d6",	x"0791",	x"07b4",	x"07bb",	
												x"07aa",	x"078f",	x"07ae",	x"078c",	
												x"07c2",	x"0783",	x"07cd",	x"0797",	
												x"07b4",	x"0794",	x"07c0",	x"079e",	
												x"07ca",	x"0771",	x"07a2",	x"0789",	
												x"0792",	x"0750",	x"07d9",	x"0786",	
												x"07d2",	x"0766",	x"07e1",	x"07b4",	
												x"07f3",	x"07aa",	x"07e1",	x"07bf",	
												x"0809",	x"07bd",	x"080c",	x"080e",	
												x"07e6",	x"07ee",	x"080d",	x"07de",	
												x"0803",	x"07e2",	x"0804",	x"07da",	
												x"07df",	x"07df",	x"0810",	x"07cb",	
												x"0835",	x"07e4",	x"0809",	x"07ea",	
												x"0816",	x"07dd",	x"0805",	x"07ed",	
												x"084b",	x"07d1",	x"084c",	x"07fa",	
												x"0818",	x"07f6",	x"07d5",	x"07de",	
												x"702f",	x"024a",	x"07f4",	x"07bf",	
												x"07ff",	x"07d8",	x"07d7",	x"07ad",	
												x"0803",	x"07bb",	x"07fc",	x"0802",	
												x"07da",	x"0777",	x"07e8",	x"07a0",	
												x"07e1",	x"07c2",	x"080c",	x"0799",	
												x"07e7",	x"07d5",	x"07e5",	x"07a9",	
												x"082b",	x"07c4",	x"07f7",	x"07e2",	
												x"0839",	x"07ec",	x"083a",	x"0810",	
												x"0855",	x"081e",	x"085b",	x"080e",	
												x"085a",	x"0856",	x"0866",	x"0816",	
												x"0852",	x"084e",	x"0856",	x"085a",	
												x"089b",	x"0843",	x"086b",	x"0859",	
												x"086c",	x"0853",	x"0886",	x"086a",	
												x"088f",	x"0825",	x"0871",	x"0884",	
												x"0899",	x"085f",	x"0893",	x"0860",	
												x"08b7",	x"086e",	x"0893",	x"0878",	
												x"05f6",	x"0887",	x"0004",	x"000a",	
												x"88b9",	x"67fa",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"124b",	
												x"0604",	x"05fe",	x"060a",	x"0618",	
												x"05f4",	x"062a",	x"05ea",	x"05eb",	
												x"05e3",	x"05e7",	x"05d5",	x"05e5",	
												x"05c0",	x"05ce",	x"05b7",	x"05d5",	
												x"05e2",	x"05da",	x"0604",	x"05fb",	
												x"0649",	x"0627",	x"0620",	x"0628",	
												x"0607",	x"0634",	x"0613",	x"062e",	
												x"060d",	x"061f",	x"05e4",	x"0639",	
												x"062f",	x"05ec",	x"0603",	x"0634",	
												x"061b",	x"0621",	x"0621",	x"0632",	
												x"0610",	x"0604",	x"0638",	x"061b",	
												x"062a",	x"0627",	x"05f8",	x"061e",	
												x"05ff",	x"0604",	x"0625",	x"060b",	
												x"0613",	x"060f",	x"062f",	x"062a",	
												x"063f",	x"0615",	x"0647",	x"062d",	
												x"0639",	x"0623",	x"0603",	x"0623",	
												x"102f",	x"124b",	x"05ea",	x"05f0",	
												x"05ec",	x"05e8",	x"05df",	x"05ef",	
												x"05d8",	x"05d8",	x"05ba",	x"05cc",	
												x"05cb",	x"05c3",	x"05d1",	x"05cf",	
												x"05c2",	x"05d9",	x"0600",	x"05cd",	
												x"0622",	x"0608",	x"0620",	x"0614",	
												x"0624",	x"062a",	x"0618",	x"0619",	
												x"0620",	x"0619",	x"05fb",	x"0615",	
												x"05d7",	x"0611",	x"0605",	x"05ee",	
												x"0600",	x"0623",	x"060f",	x"060d",	
												x"05f8",	x"0625",	x"05fb",	x"05fa",	
												x"060b",	x"0607",	x"0617",	x"0606",	
												x"05df",	x"05f8",	x"060f",	x"05fb",	
												x"0608",	x"061d",	x"060f",	x"0619",	
												x"061e",	x"061f",	x"0632",	x"0620",	
												x"063a",	x"0638",	x"0627",	x"062b",	
												x"05c2",	x"0622",	x"202f",	x"124b",	
												x"05d0",	x"05de",	x"05f5",	x"05ec",	
												x"05bb",	x"05cf",	x"05ce",	x"05dd",	
												x"05d2",	x"05d1",	x"05ac",	x"05e7",	
												x"05ae",	x"05c6",	x"05ad",	x"05bc",	
												x"05d6",	x"05dd",	x"05de",	x"05db",	
												x"0601",	x"05ea",	x"05e7",	x"05f1",	
												x"05f4",	x"05fe",	x"05fc",	x"0606",	
												x"05f7",	x"05fe",	x"05cf",	x"05df",	
												x"05ed",	x"05df",	x"05f2",	x"05e9",	
												x"0601",	x"0600",	x"0602",	x"0614",	
												x"0605",	x"05f7",	x"05f0",	x"05fb",	
												x"0617",	x"05f4",	x"05e6",	x"0600",	
												x"0607",	x"05fa",	x"0614",	x"0604",	
												x"060d",	x"0605",	x"061e",	x"05f3",	
												x"060e",	x"05fb",	x"060a",	x"060f",	
												x"0614",	x"05f4",	x"05c4",	x"0615",	
												x"302f",	x"124b",	x"05d4",	x"05a8",	
												x"05e2",	x"05d4",	x"05c7",	x"05c0",	
												x"05dd",	x"05a1",	x"05bb",	x"05c3",	
												x"05c7",	x"05a4",	x"05c6",	x"05cc",	
												x"05b0",	x"05af",	x"05e1",	x"05d1",	
												x"05e0",	x"05e7",	x"05e8",	x"05e0",	
												x"05f9",	x"05e4",	x"05f8",	x"05e7",	
												x"0604",	x"05ea",	x"05ed",	x"05ec",	
												x"05ce",	x"05eb",	x"05fb",	x"05dc",	
												x"0619",	x"0607",	x"0618",	x"0608",	
												x"0614",	x"0604",	x"060d",	x"05fd",	
												x"061b",	x"0610",	x"05ff",	x"060a",	
												x"05f0",	x"05f7",	x"061f",	x"0605",	
												x"0616",	x"0600",	x"0622",	x"05ee",	
												x"0629",	x"060d",	x"0631",	x"05fe",	
												x"0633",	x"061a",	x"0637",	x"0614",	
												x"05f4",	x"061e",	x"0004",	x"000a",	
												x"9d57",	x"caca",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"124c",	
												x"05ea",	x"05e1",	x"05f4",	x"05cf",	
												x"05e6",	x"05ef",	x"05e1",	x"05bf",	
												x"05e5",	x"05a4",	x"05d2",	x"05ca",	
												x"05d1",	x"05d0",	x"05e0",	x"05d3",	
												x"0601",	x"05a2",	x"0618",	x"0603",	
												x"0626",	x"061e",	x"061a",	x"0609",	
												x"061d",	x"0606",	x"0623",	x"061e",	
												x"0626",	x"0615",	x"061e",	x"061c",	
												x"0635",	x"0611",	x"062e",	x"062a",	
												x"0645",	x"0613",	x"0642",	x"0644",	
												x"0655",	x"063c",	x"064d",	x"064b",	
												x"0648",	x"063d",	x"0619",	x"0637",	
												x"0663",	x"0627",	x"0655",	x"064f",	
												x"066d",	x"0623",	x"0675",	x"064e",	
												x"0669",	x"064c",	x"066d",	x"064f",	
												x"0677",	x"065b",	x"05f3",	x"064b",	
												x"502f",	x"124c",	x"062a",	x"05df",	
												x"0630",	x"05f5",	x"0620",	x"05fe",	
												x"0621",	x"0600",	x"061c",	x"0603",	
												x"062b",	x"0608",	x"0633",	x"05d9",	
												x"0616",	x"05f5",	x"0650",	x"05ff",	
												x"0652",	x"0626",	x"064e",	x"0629",	
												x"065e",	x"065b",	x"064f",	x"062e",	
												x"0658",	x"0630",	x"0661",	x"063d",	
												x"0630",	x"0626",	x"0663",	x"0623",	
												x"0673",	x"065a",	x"0675",	x"0653",	
												x"0675",	x"0657",	x"0697",	x"0657",	
												x"0680",	x"065b",	x"0671",	x"064a",	
												x"0659",	x"0642",	x"0697",	x"063e",	
												x"0699",	x"0660",	x"0692",	x"0652",	
												x"0696",	x"0659",	x"0680",	x"0652",	
												x"06a1",	x"0658",	x"068c",	x"0663",	
												x"060c",	x"0650",	x"602f",	x"124c",	
												x"064c",	x"05e4",	x"0623",	x"0600",	
												x"062c",	x"05fa",	x"0634",	x"0619",	
												x"0635",	x"05f0",	x"0651",	x"05ec",	
												x"061f",	x"05fe",	x"0653",	x"05f7",	
												x"065c",	x"061c",	x"065c",	x"0638",	
												x"0666",	x"0643",	x"0668",	x"0658",	
												x"0695",	x"0652",	x"068e",	x"0669",	
												x"0695",	x"0670",	x"0664",	x"067f",	
												x"068f",	x"064d",	x"0684",	x"0682",	
												x"06a8",	x"0669",	x"069f",	x"0678",	
												x"06ac",	x"0687",	x"06a2",	x"0696",	
												x"06b9",	x"0697",	x"0687",	x"066d",	
												x"06ae",	x"068a",	x"06b2",	x"0685",	
												x"06cb",	x"0680",	x"06ba",	x"069d",	
												x"06ba",	x"0688",	x"06bc",	x"0682",	
												x"06bf",	x"0688",	x"0636",	x"0675",	
												x"702f",	x"124c",	x"065e",	x"0611",	
												x"0656",	x"063d",	x"0683",	x"0634",	
												x"069b",	x"062d",	x"067d",	x"060f",	
												x"0681",	x"063e",	x"0650",	x"0635",	
												x"0687",	x"0636",	x"068a",	x"0627",	
												x"06cd",	x"0658",	x"06e9",	x"067e",	
												x"06d7",	x"069e",	x"06d8",	x"06a3",	
												x"06c0",	x"06bc",	x"06e0",	x"06bc",	
												x"06a6",	x"06a2",	x"06f8",	x"0691",	
												x"0707",	x"06e6",	x"06fe",	x"06b0",	
												x"0708",	x"06e6",	x"0712",	x"06b9",	
												x"06f3",	x"06e6",	x"06f0",	x"06d1",	
												x"06ba",	x"06c5",	x"06ff",	x"06cc",	
												x"06f2",	x"06d3",	x"0707",	x"06df",	
												x"0733",	x"0707",	x"073b",	x"06f5",	
												x"0711",	x"06f4",	x"072f",	x"0704",	
												x"06df",	x"06fd",	x"0004",	x"000a",	
												x"d962",	x"f359",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"224d",	
												x"06db",	x"06e1",	x"06e7",	x"06b7",	
												x"06bd",	x"06c3",	x"06d3",	x"06cd",	
												x"06be",	x"06c1",	x"06d9",	x"06d8",	
												x"06ea",	x"06cd",	x"06b4",	x"06db",	
												x"06c9",	x"06bc",	x"0703",	x"06ea",	
												x"06f3",	x"0710",	x"0707",	x"0720",	
												x"0702",	x"0708",	x"0708",	x"0722",	
												x"06fe",	x"0711",	x"06d3",	x"071d",	
												x"06e0",	x"06f7",	x"0707",	x"06ea",	
												x"0715",	x"0701",	x"0704",	x"0728",	
												x"0719",	x"0706",	x"0729",	x"0711",	
												x"06ed",	x"0714",	x"06db",	x"06fc",	
												x"06f4",	x"0701",	x"0722",	x"0713",	
												x"0717",	x"070c",	x"0716",	x"0707",	
												x"0717",	x"06ef",	x"071f",	x"0706",	
												x"0710",	x"06f9",	x"06cf",	x"070a",	
												x"102f",	x"224d",	x"06c9",	x"06e2",	
												x"06be",	x"06ee",	x"06c0",	x"06b5",	
												x"069c",	x"06e8",	x"06c2",	x"0693",	
												x"06bd",	x"06bf",	x"06c4",	x"06d6",	
												x"06ad",	x"06c7",	x"06e5",	x"06c0",	
												x"06f1",	x"06e6",	x"06f1",	x"0704",	
												x"06f7",	x"0702",	x"06fe",	x"0716",	
												x"06ca",	x"06fb",	x"06d9",	x"06d8",	
												x"06c6",	x"06df",	x"06cf",	x"06c5",	
												x"06d1",	x"06d9",	x"06e5",	x"06dc",	
												x"0700",	x"06f3",	x"0716",	x"06ef",	
												x"06df",	x"0718",	x"06e9",	x"0700",	
												x"06d8",	x"0702",	x"0707",	x"070d",	
												x"0700",	x"070e",	x"06fb",	x"06f4",	
												x"0725",	x"0713",	x"0715",	x"070c",	
												x"0701",	x"071a",	x"071b",	x"0708",	
												x"0688",	x"0707",	x"202f",	x"224d",	
												x"0689",	x"06a9",	x"06be",	x"06a3",	
												x"06bd",	x"06c7",	x"069a",	x"06c3",	
												x"0691",	x"06a9",	x"06b4",	x"06af",	
												x"06b1",	x"06c6",	x"06a2",	x"06b7",	
												x"06bf",	x"06c0",	x"06e1",	x"06e8",	
												x"06e2",	x"0706",	x"06d2",	x"06e0",	
												x"06d6",	x"06e0",	x"06c9",	x"06ce",	
												x"06da",	x"06dc",	x"06ca",	x"06eb",	
												x"06e6",	x"06e8",	x"06dd",	x"06db",	
												x"06ef",	x"06d6",	x"06cb",	x"06e2",	
												x"06d5",	x"06df",	x"06f8",	x"06d0",	
												x"06f2",	x"06e0",	x"06be",	x"06db",	
												x"06e6",	x"06d6",	x"06e7",	x"06e4",	
												x"06e8",	x"06e6",	x"06e5",	x"06e5",	
												x"070d",	x"06d1",	x"06fa",	x"06f0",	
												x"06ee",	x"06e6",	x"0698",	x"06dd",	
												x"302f",	x"224d",	x"0686",	x"0669",	
												x"06a6",	x"0660",	x"0693",	x"0673",	
												x"0697",	x"067c",	x"069b",	x"0681",	
												x"06ae",	x"06a1",	x"068e",	x"06a3",	
												x"0664",	x"067f",	x"06bf",	x"0681",	
												x"06c6",	x"06ca",	x"06c2",	x"06be",	
												x"06cf",	x"06c2",	x"06d1",	x"06cd",	
												x"06de",	x"06c2",	x"06cc",	x"06bc",	
												x"069d",	x"06c3",	x"06bb",	x"06c3",	
												x"06e3",	x"06cb",	x"06db",	x"06c8",	
												x"06e5",	x"06e1",	x"06ef",	x"06ca",	
												x"06e7",	x"06d4",	x"06f8",	x"06df",	
												x"06ce",	x"06e4",	x"06f5",	x"06bb",	
												x"06e7",	x"06c4",	x"06ee",	x"06d1",	
												x"06f0",	x"06d1",	x"0713",	x"06d0",	
												x"070b",	x"06ca",	x"0707",	x"06e5",	
												x"06aa",	x"06ea",	x"0004",	x"000a",	
												x"0d65",	x"7b3a",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"224e",	
												x"06ba",	x"0684",	x"06bf",	x"06ac",	
												x"06a7",	x"0697",	x"06e5",	x"06a2",	
												x"06c7",	x"069a",	x"06c0",	x"06a0",	
												x"06ec",	x"06b6",	x"06ac",	x"06b3",	
												x"06ef",	x"06bd",	x"06fe",	x"06d1",	
												x"06ec",	x"0710",	x"06f3",	x"06fd",	
												x"06f4",	x"06e0",	x"071f",	x"06f6",	
												x"0704",	x"0701",	x"06e7",	x"06fe",	
												x"0702",	x"06d9",	x"072c",	x"06f2",	
												x"071c",	x"070f",	x"0716",	x"070a",	
												x"0725",	x"0709",	x"0721",	x"0708",	
												x"0724",	x"071d",	x"0710",	x"071e",	
												x"0739",	x"0721",	x"074a",	x"0728",	
												x"074b",	x"0725",	x"074e",	x"0741",	
												x"073e",	x"0727",	x"0739",	x"0727",	
												x"074f",	x"070f",	x"06d9",	x"072f",	
												x"502f",	x"224e",	x"070a",	x"06b1",	
												x"0724",	x"06db",	x"06ef",	x"06c9",	
												x"0700",	x"06e4",	x"0711",	x"06d8",	
												x"06fa",	x"06e6",	x"0714",	x"06cb",	
												x"06fc",	x"06e5",	x"072c",	x"06fd",	
												x"074b",	x"0708",	x"0738",	x"0725",	
												x"0720",	x"071d",	x"0750",	x"071b",	
												x"073f",	x"0741",	x"0754",	x"0701",	
												x"0724",	x"0722",	x"0740",	x"0723",	
												x"0745",	x"0718",	x"0764",	x"0729",	
												x"0748",	x"0734",	x"0761",	x"070b",	
												x"0753",	x"0735",	x"0753",	x"071d",	
												x"074e",	x"071d",	x"076c",	x"0722",	
												x"0771",	x"072a",	x"0769",	x"072f",	
												x"076e",	x"073a",	x"077d",	x"073f",	
												x"076e",	x"073b",	x"0779",	x"0739",	
												x"06f3",	x"073b",	x"602f",	x"224e",	
												x"070d",	x"06c1",	x"0710",	x"06e2",	
												x"070b",	x"0706",	x"06f9",	x"06d2",	
												x"06fb",	x"06a9",	x"0708",	x"06bc",	
												x"074e",	x"06ec",	x"0725",	x"06fb",	
												x"0757",	x"06e7",	x"0766",	x"0719",	
												x"076a",	x"0752",	x"076d",	x"0753",	
												x"0785",	x"073b",	x"07ae",	x"076a",	
												x"077f",	x"0749",	x"074d",	x"0732",	
												x"077f",	x"0723",	x"0779",	x"0751",	
												x"0782",	x"075b",	x"07a6",	x"0756",	
												x"07a5",	x"076e",	x"0785",	x"0762",	
												x"0782",	x"075b",	x"076e",	x"075d",	
												x"07a2",	x"075d",	x"07a3",	x"075b",	
												x"07a8",	x"0753",	x"07b1",	x"0768",	
												x"07b1",	x"076c",	x"07b4",	x"076d",	
												x"07a8",	x"076f",	x"075f",	x"075f",	
												x"702f",	x"224e",	x"0742",	x"06fa",	
												x"0708",	x"06f4",	x"0726",	x"06f7",	
												x"073a",	x"0718",	x"0743",	x"0717",	
												x"073d",	x"0711",	x"0737",	x"070a",	
												x"0772",	x"071e",	x"07ab",	x"0741",	
												x"077b",	x"0785",	x"07b3",	x"0771",	
												x"07b3",	x"077a",	x"07c6",	x"079d",	
												x"07cd",	x"07ad",	x"07c4",	x"077a",	
												x"077e",	x"0791",	x"07de",	x"076b",	
												x"07fc",	x"07ce",	x"0802",	x"07bb",	
												x"081c",	x"07e5",	x"0817",	x"07ce",	
												x"0808",	x"07ee",	x"0804",	x"07c7",	
												x"0801",	x"07b8",	x"0812",	x"07f0",	
												x"07fe",	x"07ed",	x"07f9",	x"07e2",	
												x"0808",	x"07e1",	x"0828",	x"0806",	
												x"0820",	x"07d5",	x"0811",	x"07fe",	
												x"06fa",	x"080c",	x"0004",	x"000a",	
												x"4bdc",	x"a570",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"324f",	
												x"06d9",	x"06f7",	x"06dd",	x"06f5",	
												x"06b8",	x"06e6",	x"06c6",	x"06b2",	
												x"06d0",	x"06b6",	x"0708",	x"06d0",	
												x"0706",	x"06e0",	x"06ba",	x"070d",	
												x"0720",	x"06d2",	x"0724",	x"0707",	
												x"0721",	x"0727",	x"06d8",	x"0730",	
												x"0703",	x"06e3",	x"070f",	x"0718",	
												x"0700",	x"0747",	x"06ed",	x"0735",	
												x"06ea",	x"0709",	x"0750",	x"0707",	
												x"0724",	x"072e",	x"0721",	x"072e",	
												x"0710",	x"070e",	x"0720",	x"071d",	
												x"070a",	x"0722",	x"0712",	x"071c",	
												x"071d",	x"0720",	x"0739",	x"072a",	
												x"070e",	x"0719",	x"0703",	x"06f5",	
												x"0711",	x"070f",	x"0734",	x"0710",	
												x"0719",	x"0727",	x"06b7",	x"070e",	
												x"102f",	x"324f",	x"06b8",	x"06cd",	
												x"06bd",	x"06d2",	x"06ac",	x"06d3",	
												x"06bf",	x"06c4",	x"06c9",	x"06c1",	
												x"06e0",	x"06d7",	x"06df",	x"06e6",	
												x"06b7",	x"06d9",	x"0719",	x"06df",	
												x"070e",	x"071d",	x"06f0",	x"0704",	
												x"0707",	x"06f1",	x"06f9",	x"0702",	
												x"070e",	x"071d",	x"06ff",	x"0704",	
												x"06db",	x"0703",	x"06e3",	x"0700",	
												x"070b",	x"0702",	x"06f8",	x"072a",	
												x"06f7",	x"0706",	x"06f6",	x"06f9",	
												x"06f4",	x"0733",	x"06eb",	x"0719",	
												x"06cd",	x"06fa",	x"06f9",	x"06e8",	
												x"0710",	x"0704",	x"0712",	x"0704",	
												x"071d",	x"071a",	x"0713",	x"0704",	
												x"0717",	x"0717",	x"072f",	x"0728",	
												x"06ab",	x"0727",	x"202f",	x"324f",	
												x"06aa",	x"06bc",	x"06b1",	x"06bd",	
												x"06b7",	x"069d",	x"06c6",	x"06c0",	
												x"06c7",	x"06da",	x"06d3",	x"0700",	
												x"06c7",	x"06ef",	x"06b3",	x"06e2",	
												x"06d1",	x"06eb",	x"06e7",	x"0714",	
												x"06f0",	x"0702",	x"06d8",	x"0704",	
												x"06ec",	x"06e1",	x"06ce",	x"06f2",	
												x"0700",	x"06db",	x"06c3",	x"06e8",	
												x"06e7",	x"06dc",	x"06fc",	x"06e7",	
												x"06f8",	x"06f0",	x"06dd",	x"06f0",	
												x"06ee",	x"06d6",	x"06fe",	x"06fd",	
												x"0705",	x"06f5",	x"06d5",	x"06ee",	
												x"0709",	x"06fb",	x"06fd",	x"06f7",	
												x"0708",	x"06e8",	x"06e5",	x"06f9",	
												x"0702",	x"06e4",	x"0704",	x"06fe",	
												x"0720",	x"06e8",	x"0684",	x"06ec",	
												x"302f",	x"324f",	x"068b",	x"0675",	
												x"068d",	x"067f",	x"0680",	x"0675",	
												x"06a1",	x"069c",	x"06a6",	x"0685",	
												x"06ab",	x"06a3",	x"06b5",	x"0688",	
												x"0696",	x"06cd",	x"06d5",	x"06b4",	
												x"06c3",	x"06c7",	x"06d8",	x"06c9",	
												x"06df",	x"06c0",	x"06dd",	x"06e0",	
												x"06d3",	x"06d6",	x"06c5",	x"06da",	
												x"06a6",	x"06ce",	x"06e2",	x"06df",	
												x"06eb",	x"06cd",	x"06e8",	x"06cc",	
												x"06fe",	x"06f3",	x"0704",	x"06de",	
												x"06fb",	x"06f2",	x"06f8",	x"06f7",	
												x"06f4",	x"06e8",	x"071a",	x"070a",	
												x"0701",	x"070e",	x"06fd",	x"06e6",	
												x"0712",	x"06e8",	x"0701",	x"06f1",	
												x"0702",	x"06db",	x"070f",	x"06e7",	
												x"06cb",	x"06eb",	x"0004",	x"000a",	
												x"14a8",	x"c453",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"3250",	
												x"06c1",	x"0689",	x"06b5",	x"06aa",	
												x"06be",	x"068a",	x"06a6",	x"06c1",	
												x"06be",	x"069f",	x"06c7",	x"06c7",	
												x"06ca",	x"06c6",	x"06cc",	x"06f0",	
												x"0707",	x"06dd",	x"070c",	x"06eb",	
												x"0717",	x"06fb",	x"0704",	x"0707",	
												x"070e",	x"06fa",	x"071f",	x"06fb",	
												x"0720",	x"0713",	x"06f1",	x"0711",	
												x"072a",	x"06fe",	x"0720",	x"0709",	
												x"0731",	x"073a",	x"072e",	x"071e",	
												x"072c",	x"0719",	x"0728",	x"071f",	
												x"074b",	x"071e",	x"0724",	x"071a",	
												x"0775",	x"073d",	x"0745",	x"0730",	
												x"074e",	x"072c",	x"0734",	x"0730",	
												x"0752",	x"0715",	x"0763",	x"071b",	
												x"0767",	x"0741",	x"06e5",	x"0719",	
												x"502f",	x"3250",	x"0704",	x"06e8",	
												x"06fa",	x"06d7",	x"06fe",	x"06c3",	
												x"0714",	x"06c4",	x"0711",	x"06cd",	
												x"0704",	x"0705",	x"0733",	x"06f3",	
												x"070f",	x"072a",	x"0736",	x"0723",	
												x"0755",	x"0720",	x"0751",	x"0750",	
												x"0740",	x"0748",	x"0745",	x"072a",	
												x"0745",	x"072f",	x"0748",	x"0739",	
												x"0728",	x"071a",	x"076a",	x"0725",	
												x"076d",	x"0744",	x"0753",	x"0738",	
												x"0752",	x"0728",	x"0766",	x"072b",	
												x"0778",	x"073d",	x"07a6",	x"0739",	
												x"0752",	x"0747",	x"079b",	x"0741",	
												x"076f",	x"074d",	x"0776",	x"074e",	
												x"0781",	x"074b",	x"07a3",	x"0754",	
												x"077e",	x"075f",	x"07ad",	x"0760",	
												x"06fd",	x"074d",	x"602f",	x"3250",	
												x"072c",	x"06db",	x"071f",	x"06e8",	
												x"06e9",	x"06d2",	x"072c",	x"06dc",	
												x"0723",	x"06ea",	x"071b",	x"06ff",	
												x"072d",	x"06f0",	x"0726",	x"071d",	
												x"0776",	x"0711",	x"0789",	x"0737",	
												x"0778",	x"073b",	x"078f",	x"0745",	
												x"0780",	x"072b",	x"077e",	x"0759",	
												x"077e",	x"0751",	x"076c",	x"0784",	
												x"0782",	x"0746",	x"078f",	x"0760",	
												x"0794",	x"076b",	x"0794",	x"0756",	
												x"0784",	x"0757",	x"07a3",	x"077e",	
												x"07b3",	x"076c",	x"0781",	x"0771",	
												x"0792",	x"0774",	x"07b5",	x"077e",	
												x"07ba",	x"0781",	x"07b1",	x"078a",	
												x"07e3",	x"077b",	x"07e1",	x"0790",	
												x"07e2",	x"078f",	x"073a",	x"0771",	
												x"702f",	x"3250",	x"0738",	x"0705",	
												x"0736",	x"0716",	x"0745",	x"0701",	
												x"0786",	x"0703",	x"0752",	x"0717",	
												x"074f",	x"0726",	x"0756",	x"0716",	
												x"0759",	x"073b",	x"07af",	x"073e",	
												x"07b5",	x"0778",	x"07c2",	x"077b",	
												x"07b2",	x"07b0",	x"07cf",	x"0799",	
												x"07d4",	x"077e",	x"07e4",	x"07a3",	
												x"07b5",	x"077e",	x"07ea",	x"078a",	
												x"07ec",	x"07b0",	x"0807",	x"07a4",	
												x"0832",	x"07e3",	x"07fd",	x"07cf",	
												x"0802",	x"07f2",	x"081c",	x"07f2",	
												x"07e6",	x"07dc",	x"0820",	x"07ea",	
												x"0818",	x"07fa",	x"0817",	x"080a",	
												x"083d",	x"07e1",	x"0839",	x"0808",	
												x"0847",	x"07fe",	x"0827",	x"07fd",	
												x"0603",	x"07ef",	x"0004",	x"000a",	
												x"5225",	x"ed43",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"0251",	
												x"08c0",	x"06f6",	x"07ca",	x"06c9",	
												x"0503",	x"07b2",	x"062f",	x"03e7",	
												x"079c",	x"05ae",	x"0692",	x"08c8",	
												x"071d",	x"0839",	x"0482",	x"076e",	
												x"0883",	x"0718",	x"052f",	x"0861",	
												x"045f",	x"08cc",	x"0855",	x"0895",	
												x"0894",	x"07d7",	x"0691",	x"08fc",	
												x"08a1",	x"07b6",	x"059d",	x"0504",	
												x"0592",	x"06d5",	x"0583",	x"03a4",	
												x"0882",	x"067d",	x"0575",	x"0707",	
												x"0704",	x"04d7",	x"070f",	x"07e2",	
												x"06c8",	x"0892",	x"056a",	x"07b5",	
												x"082b",	x"0518",	x"072d",	x"061a",	
												x"0846",	x"060c",	x"068d",	x"0943",	
												x"06b2",	x"064f",	x"07e9",	x"05cc",	
												x"02fc",	x"05fa",	x"06e0",	x"063f",	
												x"1030",	x"0251",	x"069b",	x"08a9",	
												x"0732",	x"06af",	x"07fd",	x"06c6",	
												x"05d9",	x"08c2",	x"053c",	x"05a3",	
												x"0477",	x"07ba",	x"08cc",	x"0823",	
												x"0325",	x"06e3",	x"05e1",	x"04d8",	
												x"061f",	x"0584",	x"05bf",	x"0865",	
												x"0687",	x"074d",	x"07dd",	x"0748",	
												x"0433",	x"06ca",	x"05b1",	x"0566",	
												x"085b",	x"05b5",	x"062f",	x"080e",	
												x"0652",	x"0676",	x"075f",	x"06d1",	
												x"06e9",	x"0628",	x"03cd",	x"0764",	
												x"05a8",	x"05de",	x"0747",	x"06df",	
												x"04df",	x"05bf",	x"048d",	x"0705",	
												x"06b8",	x"064d",	x"0651",	x"068d",	
												x"0818",	x"0849",	x"0679",	x"05ee",	
												x"075f",	x"0650",	x"0861",	x"082b",	
												x"07dc",	x"04ec",	x"2030",	x"0251",	
												x"07be",	x"0480",	x"07cb",	x"07dc",	
												x"07dd",	x"07ea",	x"07d4",	x"082e",	
												x"07cd",	x"080a",	x"07c2",	x"07d4",	
												x"07be",	x"07d4",	x"0805",	x"0815",	
												x"07fe",	x"0813",	x"07c8",	x"081e",	
												x"07a9",	x"07aa",	x"07a7",	x"07b0",	
												x"0790",	x"07ae",	x"07c2",	x"07b5",	
												x"07c3",	x"076e",	x"07e8",	x"07f0",	
												x"07a7",	x"058d",	x"07ad",	x"0790",	
												x"07c1",	x"076f",	x"0755",	x"07c8",	
												x"06b5",	x"0774",	x"07a8",	x"0764",	
												x"0712",	x"0787",	x"07cf",	x"075e",	
												x"0555",	x"06d5",	x"070f",	x"0730",	
												x"059f",	x"07d9",	x"07f2",	x"078a",	
												x"07e0",	x"0825",	x"07bf",	x"07dd",	
												x"0822",	x"07e3",	x"07d7",	x"0800",	
												x"3030",	x"0251",	x"07aa",	x"07c0",	
												x"07ff",	x"07de",	x"07d2",	x"07ea",	
												x"07d2",	x"07c1",	x"07c8",	x"07cc",	
												x"07de",	x"07aa",	x"07d6",	x"07e3",	
												x"07ec",	x"07df",	x"079c",	x"07d8",	
												x"07ae",	x"07b5",	x"078d",	x"07aa",	
												x"07a3",	x"07c2",	x"0783",	x"0798",	
												x"07a5",	x"07a6",	x"07bc",	x"07c6",	
												x"07f2",	x"07ba",	x"0746",	x"079c",	
												x"07b8",	x"0793",	x"07ba",	x"0792",	
												x"0775",	x"0780",	x"0777",	x"07ae",	
												x"0786",	x"076b",	x"078d",	x"0797",	
												x"07d7",	x"07c3",	x"07bd",	x"07ac",	
												x"07c6",	x"0790",	x"07d5",	x"07c7",	
												x"07e0",	x"07e2",	x"0803",	x"07e2",	
												x"07fa",	x"07e7",	x"0800",	x"07d2",	
												x"07bf",	x"07e9",	x"0004",	x"000a",	
												x"2c0c",	x"2d73",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"0252",	
												x"07de",	x"07a6",	x"07ee",	x"07d6",	
												x"07e5",	x"07e6",	x"07f8",	x"07e3",	
												x"07e9",	x"0813",	x"07f6",	x"07ed",	
												x"07f7",	x"07f4",	x"0824",	x"080a",	
												x"07ce",	x"082b",	x"07c2",	x"07e2",	
												x"07a2",	x"07d9",	x"07c7",	x"07c9",	
												x"07dd",	x"07d5",	x"07c9",	x"07d2",	
												x"07f4",	x"07c9",	x"0804",	x"0807",	
												x"07dd",	x"07e4",	x"07e2",	x"07e1",	
												x"07ee",	x"07d5",	x"07e9",	x"07b8",	
												x"07d7",	x"07f5",	x"07e6",	x"07ca",	
												x"07e0",	x"07dd",	x"0819",	x"07f5",	
												x"0804",	x"0801",	x"07fe",	x"07ff",	
												x"07f5",	x"07fd",	x"082a",	x"0812",	
												x"0842",	x"081f",	x"0836",	x"0831",	
												x"085e",	x"0827",	x"0828",	x"083c",	
												x"5030",	x"0252",	x"083c",	x"07f3",	
												x"0863",	x"083a",	x"0862",	x"0856",	
												x"0840",	x"0852",	x"083d",	x"083f",	
												x"085b",	x"085a",	x"0844",	x"085e",	
												x"0858",	x"085f",	x"082f",	x"0834",	
												x"0823",	x"0817",	x"0804",	x"081e",	
												x"0801",	x"080b",	x"0806",	x"0807",	
												x"080b",	x"0801",	x"0835",	x"0803",	
												x"0824",	x"0833",	x"081e",	x"0808",	
												x"07ea",	x"080f",	x"07e9",	x"07c7",	
												x"07fc",	x"07e3",	x"0805",	x"07e4",	
												x"081b",	x"07d6",	x"085c",	x"07ef",	
												x"0855",	x"0839",	x"0854",	x"083e",	
												x"084b",	x"0828",	x"084c",	x"0823",	
												x"086f",	x"0800",	x"0883",	x"083f",	
												x"089c",	x"084f",	x"0897",	x"085f",	
												x"0844",	x"0868",	x"6030",	x"0252",	
												x"084e",	x"0808",	x"0864",	x"0866",	
												x"0868",	x"0860",	x"0870",	x"085c",	
												x"0871",	x"085f",	x"0879",	x"086b",	
												x"085e",	x"0864",	x"087c",	x"085e",	
												x"0845",	x"0840",	x"083d",	x"0856",	
												x"0838",	x"0840",	x"0843",	x"082f",	
												x"0828",	x"07f3",	x"0844",	x"0819",	
												x"0856",	x"081e",	x"0885",	x"0852",	
												x"0843",	x"0865",	x"0852",	x"084a",	
												x"0848",	x"083a",	x"085c",	x"083d",	
												x"0839",	x"0814",	x"0859",	x"0843",	
												x"086a",	x"0849",	x"08a4",	x"082c",	
												x"08af",	x"0871",	x"087b",	x"0856",	
												x"0891",	x"0846",	x"08b5",	x"0855",	
												x"08be",	x"087e",	x"08d1",	x"08af",	
												x"08d7",	x"0891",	x"08c7",	x"088f",	
												x"7030",	x"0252",	x"08bc",	x"0871",	
												x"08f5",	x"08c4",	x"08b6",	x"08ce",	
												x"08cf",	x"08da",	x"08dd",	x"08e0",	
												x"08ce",	x"08e2",	x"08b5",	x"08da",	
												x"08ff",	x"08cf",	x"08c0",	x"08dd",	
												x"08aa",	x"08d7",	x"08b8",	x"08aa",	
												x"08bb",	x"08a9",	x"08b3",	x"089f",	
												x"08ac",	x"08b6",	x"08b0",	x"08ad",	
												x"08da",	x"08dc",	x"087c",	x"08bb",	
												x"08d4",	x"0896",	x"0908",	x"089f",	
												x"08c6",	x"08c4",	x"08bc",	x"08a0",	
												x"0913",	x"08b8",	x"08bd",	x"08dc",	
												x"0913",	x"08cc",	x"08fc",	x"0914",	
												x"093d",	x"08e8",	x"0933",	x"091a",	
												x"0958",	x"08f2",	x"0966",	x"0917",	
												x"0961",	x"094a",	x"0953",	x"0956",	
												x"05c2",	x"093f",	x"0004",	x"000a",	
												x"cd49",	x"b45b",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"1253",	
												x"05ce",	x"05cd",	x"05e0",	x"05dd",	
												x"05f0",	x"0608",	x"05fc",	x"05fb",	
												x"05ec",	x"05ec",	x"05ff",	x"05f5",	
												x"0611",	x"0611",	x"05cc",	x"0615",	
												x"060c",	x"060b",	x"061c",	x"0618",	
												x"061a",	x"0610",	x"05f9",	x"0629",	
												x"05f9",	x"061a",	x"05fb",	x"0606",	
												x"05ff",	x"0614",	x"05de",	x"0609",	
												x"0602",	x"05e9",	x"0606",	x"0621",	
												x"0605",	x"060d",	x"0609",	x"0603",	
												x"0607",	x"0606",	x"0609",	x"0610",	
												x"060a",	x"05f4",	x"05d8",	x"0622",	
												x"060f",	x"05e6",	x"061c",	x"0608",	
												x"061e",	x"062d",	x"063c",	x"0621",	
												x"0639",	x"061c",	x"0632",	x"0638",	
												x"0636",	x"05fa",	x"05db",	x"0620",	
												x"1030",	x"1253",	x"05cd",	x"05f3",	
												x"05ce",	x"05da",	x"05dc",	x"05d1",	
												x"05ee",	x"05d1",	x"05ee",	x"05fd",	
												x"05fa",	x"05f1",	x"0613",	x"0616",	
												x"05df",	x"0624",	x"05f8",	x"05ef",	
												x"060d",	x"0613",	x"060f",	x"060c",	
												x"0617",	x"0612",	x"060e",	x"061c",	
												x"0605",	x"061c",	x"0601",	x"060d",	
												x"05d1",	x"05e2",	x"05e0",	x"05ed",	
												x"05fa",	x"0604",	x"0607",	x"0612",	
												x"05f7",	x"0622",	x"05f8",	x"0609",	
												x"0619",	x"05fb",	x"0611",	x"0617",	
												x"05e2",	x"0606",	x"062f",	x"0604",	
												x"061c",	x"062a",	x"062a",	x"062d",	
												x"061e",	x"0632",	x"0629",	x"060b",	
												x"0628",	x"0636",	x"0621",	x"0616",	
												x"05c1",	x"062f",	x"2030",	x"1253",	
												x"05bd",	x"05c3",	x"05da",	x"05d0",	
												x"05d2",	x"05c6",	x"05ca",	x"05d3",	
												x"05bd",	x"05bc",	x"05fb",	x"0605",	
												x"0607",	x"0605",	x"05e7",	x"0605",	
												x"05f1",	x"0601",	x"05fa",	x"060b",	
												x"0605",	x"061a",	x"05f4",	x"05fc",	
												x"05e3",	x"0606",	x"05e9",	x"05e4",	
												x"05dd",	x"05eb",	x"05b7",	x"05ec",	
												x"05ef",	x"05ce",	x"05ff",	x"05f1",	
												x"060b",	x"05fb",	x"0607",	x"060f",	
												x"0604",	x"05f9",	x"05fe",	x"060d",	
												x"0609",	x"0602",	x"05da",	x"05ff",	
												x"05ff",	x"05b6",	x"060d",	x"05f7",	
												x"060c",	x"05fd",	x"0619",	x"0602",	
												x"0616",	x"0608",	x"0605",	x"0616",	
												x"0619",	x"05fb",	x"05b4",	x"05f9",	
												x"3030",	x"1253",	x"05ba",	x"05eb",	
												x"05c4",	x"05a3",	x"05d4",	x"05c2",	
												x"05e6",	x"05d3",	x"05e3",	x"05dd",	
												x"05cb",	x"05f2",	x"05f1",	x"05e0",	
												x"05b4",	x"05ef",	x"05de",	x"05e4",	
												x"05f8",	x"05df",	x"05f4",	x"05ff",	
												x"05f2",	x"05e8",	x"05e2",	x"05ec",	
												x"0600",	x"05f0",	x"05d6",	x"05e7",	
												x"05ac",	x"05b8",	x"05ec",	x"05c6",	
												x"05f9",	x"05fe",	x"0607",	x"05f9",	
												x"0612",	x"05fe",	x"05f2",	x"0600",	
												x"05f8",	x"05fe",	x"05fe",	x"05d2",	
												x"05f1",	x"05fc",	x"0617",	x"05dc",	
												x"0605",	x"0605",	x"0610",	x"0600",	
												x"0619",	x"05f8",	x"062f",	x"0601",	
												x"062f",	x"0614",	x"062b",	x"0612",	
												x"05db",	x"05fb",	x"0004",	x"000a",	
												x"9c4a",	x"cb7e",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"1254",	
												x"05e0",	x"05d5",	x"0602",	x"05e1",	
												x"05ec",	x"05de",	x"0607",	x"05df",	
												x"0603",	x"05dc",	x"05e6",	x"05ff",	
												x"05f5",	x"05e6",	x"0600",	x"05fc",	
												x"05ff",	x"05fd",	x"0609",	x"061a",	
												x"0604",	x"0621",	x"0605",	x"0609",	
												x"060a",	x"05fe",	x"0605",	x"0619",	
												x"05fe",	x"0608",	x"05f6",	x"060f",	
												x"061d",	x"060f",	x"0635",	x"060a",	
												x"0643",	x"063a",	x"064f",	x"0641",	
												x"063c",	x"0635",	x"062f",	x"062f",	
												x"062b",	x"0623",	x"061e",	x"0624",	
												x"0627",	x"061c",	x"064f",	x"0629",	
												x"064f",	x"063d",	x"0659",	x"065a",	
												x"0655",	x"0649",	x"064d",	x"0640",	
												x"066f",	x"065c",	x"0608",	x"065b",	
												x"5030",	x"1254",	x"061b",	x"05f5",	
												x"0636",	x"0600",	x"0621",	x"05eb",	
												x"062f",	x"0617",	x"0638",	x"062a",	
												x"0636",	x"0623",	x"0635",	x"063b",	
												x"0639",	x"064b",	x"064a",	x"061d",	
												x"0656",	x"064a",	x"064a",	x"064c",	
												x"065f",	x"064a",	x"065a",	x"064a",	
												x"0656",	x"0653",	x"0644",	x"0634",	
												x"063d",	x"0632",	x"064f",	x"062d",	
												x"0657",	x"0648",	x"0652",	x"0655",	
												x"065e",	x"0649",	x"066a",	x"0655",	
												x"067b",	x"0657",	x"0677",	x"063a",	
												x"0659",	x"0651",	x"0659",	x"063f",	
												x"0688",	x"065d",	x"0671",	x"0655",	
												x"0698",	x"065c",	x"0689",	x"0663",	
												x"0688",	x"0685",	x"0678",	x"065d",	
												x"063f",	x"0655",	x"6030",	x"1254",	
												x"062b",	x"0608",	x"0632",	x"0614",	
												x"062e",	x"0608",	x"0642",	x"060e",	
												x"0647",	x"0636",	x"0665",	x"062d",	
												x"0662",	x"0648",	x"065e",	x"0651",	
												x"066b",	x"064f",	x"0679",	x"0657",	
												x"0664",	x"0651",	x"067a",	x"0668",	
												x"067b",	x"066a",	x"0664",	x"066b",	
												x"0686",	x"065c",	x"0671",	x"066b",	
												x"067e",	x"064b",	x"0676",	x"0667",	
												x"0694",	x"0671",	x"069e",	x"0688",	
												x"06aa",	x"0683",	x"0694",	x"0672",	
												x"06a0",	x"0680",	x"0687",	x"0691",	
												x"0687",	x"0680",	x"068f",	x"067d",	
												x"06ba",	x"067e",	x"06b5",	x"0696",	
												x"06b9",	x"068e",	x"06ae",	x"068c",	
												x"06b6",	x"0695",	x"067d",	x"0683",	
												x"7030",	x"1254",	x"068c",	x"0642",	
												x"0679",	x"065b",	x"067f",	x"0633",	
												x"06b3",	x"067b",	x"06bb",	x"0676",	
												x"06bb",	x"068b",	x"06b3",	x"068e",	
												x"06a1",	x"06a1",	x"06cd",	x"0684",	
												x"06d5",	x"06c8",	x"06d1",	x"06be",	
												x"06c8",	x"06cc",	x"06d9",	x"06bc",	
												x"06d2",	x"06d2",	x"06bf",	x"06bb",	
												x"06a5",	x"06cc",	x"06f6",	x"06c4",	
												x"0704",	x"06db",	x"06f9",	x"06dc",	
												x"06f1",	x"06e2",	x"0707",	x"06f3",	
												x"06f7",	x"06f8",	x"06f9",	x"0701",	
												x"06c7",	x"06f6",	x"06fd",	x"06d9",	
												x"070c",	x"06eb",	x"070d",	x"06e8",	
												x"073f",	x"0718",	x"0745",	x"0715",	
												x"0744",	x"0736",	x"0720",	x"0707",	
												x"06c5",	x"0716",	x"0004",	x"000a",	
												x"d911",	x"fd22",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"2255",	
												x"06af",	x"06ec",	x"06cb",	x"06c7",	
												x"06cb",	x"06c3",	x"06d9",	x"06de",	
												x"06e1",	x"06e3",	x"0727",	x"06ff",	
												x"06f2",	x"0737",	x"06c5",	x"06f0",	
												x"070a",	x"06c9",	x"070c",	x"071c",	
												x"06e2",	x"06f8",	x"071e",	x"071d",	
												x"06d9",	x"0703",	x"06ef",	x"06fe",	
												x"06fe",	x"070f",	x"06b5",	x"06ff",	
												x"06dc",	x"06e3",	x"06f5",	x"0704",	
												x"06df",	x"06ee",	x"06e6",	x"06f8",	
												x"0719",	x"0715",	x"0708",	x"0716",	
												x"0705",	x"0702",	x"06c6",	x"06ef",	
												x"06ec",	x"06da",	x"06f5",	x"0707",	
												x"06ee",	x"06f8",	x"072e",	x"06fb",	
												x"0721",	x"0708",	x"070d",	x"0702",	
												x"072b",	x"0707",	x"0699",	x"0703",	
												x"1030",	x"2255",	x"06aa",	x"06ab",	
												x"06dc",	x"06c0",	x"06ae",	x"06db",	
												x"06a3",	x"06ca",	x"06b6",	x"06c9",	
												x"06e8",	x"06d9",	x"06f1",	x"0706",	
												x"06a9",	x"06f1",	x"06f9",	x"06ec",	
												x"06f5",	x"06f3",	x"06ed",	x"06ee",	
												x"06f4",	x"06fa",	x"06f5",	x"06f1",	
												x"06d1",	x"06fd",	x"06ca",	x"06e0",	
												x"06c1",	x"06ec",	x"06e4",	x"06bc",	
												x"06f4",	x"06f6",	x"06ee",	x"0711",	
												x"06d2",	x"0703",	x"0716",	x"06ec",	
												x"070c",	x"0706",	x"06e7",	x"0705",	
												x"06a6",	x"06e0",	x"06f6",	x"06e5",	
												x"06db",	x"06eb",	x"06fe",	x"06e0",	
												x"071a",	x"06f2",	x"072f",	x"0714",	
												x"06f5",	x"0724",	x"0723",	x"06fe",	
												x"06be",	x"0715",	x"2030",	x"2255",	
												x"06a8",	x"06c9",	x"067d",	x"06a7",	
												x"06a2",	x"06b5",	x"06a8",	x"06bb",	
												x"06a1",	x"06b1",	x"06cc",	x"06d6",	
												x"06c2",	x"06ce",	x"067f",	x"06d4",	
												x"06d9",	x"06d3",	x"06d2",	x"06f1",	
												x"06d0",	x"06e9",	x"06c8",	x"06df",	
												x"06d4",	x"06df",	x"06c4",	x"06f8",	
												x"06c8",	x"06bb",	x"0671",	x"06dc",	
												x"06bd",	x"06b7",	x"06cb",	x"06ba",	
												x"06cd",	x"06c8",	x"06c1",	x"06cb",	
												x"06fa",	x"0696",	x"06f4",	x"06ec",	
												x"06ef",	x"06dc",	x"06c5",	x"06d0",	
												x"06d7",	x"06c7",	x"06d4",	x"06dd",	
												x"06e2",	x"06da",	x"06e0",	x"06ea",	
												x"06e5",	x"06db",	x"06f8",	x"06d2",	
												x"06f2",	x"06e4",	x"066b",	x"06dd",	
												x"3030",	x"2255",	x"069b",	x"068c",	
												x"0698",	x"069f",	x"0693",	x"0687",	
												x"069e",	x"0690",	x"06b2",	x"069c",	
												x"06b3",	x"06b4",	x"0688",	x"06ce",	
												x"0676",	x"06ac",	x"06b7",	x"06b7",	
												x"06d2",	x"06d2",	x"06d0",	x"06c8",	
												x"06d5",	x"06b8",	x"06ca",	x"06c2",	
												x"06c6",	x"06bc",	x"06ac",	x"06b2",	
												x"0691",	x"06b0",	x"06a5",	x"06a8",	
												x"06c2",	x"06c1",	x"06c4",	x"06af",	
												x"06cb",	x"06ca",	x"06d9",	x"06b7",	
												x"06d6",	x"06e5",	x"06eb",	x"06db",	
												x"06b7",	x"06cc",	x"06fd",	x"06c2",	
												x"06ce",	x"06cf",	x"06fa",	x"06cf",	
												x"06f9",	x"06ec",	x"070d",	x"06d6",	
												x"06fc",	x"06be",	x"06f9",	x"06ce",	
												x"0685",	x"06df",	x"0004",	x"000a",	
												x"0abd",	x"7be0",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"2256",	
												x"0678",	x"0695",	x"06c8",	x"068a",	
												x"06b4",	x"06b9",	x"06c4",	x"06ba",	
												x"06b4",	x"06b3",	x"06c1",	x"06a2",	
												x"06c9",	x"06d9",	x"06d2",	x"06d3",	
												x"06e6",	x"06d9",	x"06e3",	x"06e0",	
												x"06de",	x"06f4",	x"06f5",	x"06ed",	
												x"06cd",	x"06f2",	x"06f7",	x"06f0",	
												x"06ee",	x"06ef",	x"06e9",	x"06f5",	
												x"06fe",	x"06f7",	x"06ff",	x"071f",	
												x"0703",	x"0715",	x"06f5",	x"0702",	
												x"0703",	x"06fb",	x"0715",	x"06f5",	
												x"0709",	x"0709",	x"0703",	x"0705",	
												x"0712",	x"0706",	x"0717",	x"0708",	
												x"071e",	x"0711",	x"072e",	x"0719",	
												x"0722",	x"0712",	x"0737",	x"0717",	
												x"073f",	x"071b",	x"06d7",	x"0734",	
												x"5030",	x"2256",	x"06fa",	x"06e5",	
												x"06ea",	x"06f3",	x"06de",	x"06fc",	
												x"070c",	x"06bf",	x"06e6",	x"06dc",	
												x"06fb",	x"06e5",	x"0715",	x"06fd",	
												x"0709",	x"070e",	x"071a",	x"0713",	
												x"0736",	x"072c",	x"0720",	x"072e",	
												x"0711",	x"071f",	x"070b",	x"0720",	
												x"0711",	x"0714",	x"0710",	x"0713",	
												x"06ee",	x"06f8",	x"0720",	x"06dc",	
												x"072e",	x"0720",	x"0746",	x"0711",	
												x"0737",	x"073c",	x"0739",	x"070a",	
												x"074e",	x"0724",	x"0731",	x"072c",	
												x"0731",	x"071e",	x"0764",	x"0729",	
												x"0756",	x"0733",	x"0751",	x"072e",	
												x"077f",	x"073c",	x"0772",	x"073d",	
												x"075e",	x"0741",	x"075f",	x"0744",	
												x"06e4",	x"074a",	x"6030",	x"2256",	
												x"06fc",	x"06d8",	x"0703",	x"06f1",	
												x"0707",	x"06ea",	x"0737",	x"06f1",	
												x"0714",	x"070a",	x"071e",	x"0706",	
												x"0723",	x"0713",	x"0739",	x"072e",	
												x"0756",	x"0733",	x"0760",	x"0750",	
												x"0733",	x"0752",	x"0750",	x"0743",	
												x"0754",	x"0751",	x"0767",	x"0748",	
												x"0766",	x"0735",	x"0747",	x"0741",	
												x"0741",	x"0737",	x"0777",	x"0757",	
												x"0784",	x"076f",	x"076e",	x"076e",	
												x"0781",	x"0763",	x"078c",	x"075b",	
												x"0788",	x"077a",	x"0771",	x"077b",	
												x"0783",	x"076d",	x"078f",	x"076a",	
												x"0796",	x"075d",	x"07b8",	x"077a",	
												x"07aa",	x"0779",	x"07b1",	x"077b",	
												x"07b7",	x"078f",	x"0721",	x"077d",	
												x"7030",	x"2256",	x"0765",	x"0738",	
												x"072d",	x"0732",	x"0770",	x"0728",	
												x"0788",	x"075a",	x"07a5",	x"0770",	
												x"0791",	x"079b",	x"077e",	x"078a",	
												x"0778",	x"0783",	x"07b7",	x"0778",	
												x"07d3",	x"07d3",	x"07b3",	x"07cd",	
												x"07ba",	x"07b8",	x"07b1",	x"07c3",	
												x"07d9",	x"07a9",	x"07bc",	x"07c5",	
												x"07b1",	x"07bf",	x"07ca",	x"07b6",	
												x"07fe",	x"07d9",	x"07f7",	x"07db",	
												x"080c",	x"07ff",	x"07fb",	x"07e4",	
												x"07f4",	x"0803",	x"07e1",	x"07e7",	
												x"07e0",	x"07cf",	x"07f4",	x"07ea",	
												x"0821",	x"07f3",	x"080e",	x"07f3",	
												x"0840",	x"0801",	x"083b",	x"0809",	
												x"084b",	x"0844",	x"0819",	x"081f",	
												x"06ce",	x"0832",	x"0004",	x"000a",	
												x"46ef",	x"aef4",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"3257",	
												x"06b2",	x"06f8",	x"06de",	x"06d0",	
												x"06b1",	x"06d0",	x"06b2",	x"06c7",	
												x"06a9",	x"06d2",	x"06f1",	x"06cd",	
												x"06f0",	x"06e8",	x"06e6",	x"0710",	
												x"06d8",	x"0714",	x"0702",	x"070b",	
												x"06f9",	x"070f",	x"06f1",	x"071b",	
												x"0720",	x"0707",	x"06f8",	x"070d",	
												x"0710",	x"0704",	x"06c1",	x"072a",	
												x"06ee",	x"06df",	x"0710",	x"0708",	
												x"06f3",	x"06fb",	x"06f7",	x"0706",	
												x"0703",	x"06fc",	x"0709",	x"06e4",	
												x"070e",	x"0707",	x"06e6",	x"06fc",	
												x"06f6",	x"06ed",	x"0709",	x"0718",	
												x"06eb",	x"06f6",	x"06fd",	x"06d2",	
												x"0707",	x"0707",	x"0735",	x"070b",	
												x"06f7",	x"0728",	x"06b0",	x"06fa",	
												x"1030",	x"3257",	x"067a",	x"06ae",	
												x"06a2",	x"06a4",	x"067f",	x"06be",	
												x"06be",	x"06cb",	x"06b3",	x"06dc",	
												x"06eb",	x"06d4",	x"06f9",	x"06dd",	
												x"06c3",	x"06f5",	x"06fb",	x"06d7",	
												x"06e1",	x"0705",	x"06bf",	x"06e8",	
												x"0734",	x"06dc",	x"06d3",	x"0705",	
												x"06ee",	x"06ef",	x"06d9",	x"06e8",	
												x"06ba",	x"06ee",	x"06d5",	x"06ef",	
												x"06dc",	x"06f7",	x"06e5",	x"06e0",	
												x"06e7",	x"06e7",	x"06d2",	x"06f7",	
												x"06e2",	x"06f9",	x"06ef",	x"06fa",	
												x"06e1",	x"06f6",	x"06f1",	x"06d4",	
												x"06f4",	x"06eb",	x"06f2",	x"06e0",	
												x"06fc",	x"06f9",	x"071a",	x"06fb",	
												x"0728",	x"0721",	x"071a",	x"072c",	
												x"06b8",	x"0712",	x"2030",	x"3257",	
												x"069d",	x"06df",	x"06a3",	x"06b2",	
												x"06ad",	x"06b1",	x"06aa",	x"06b5",	
												x"06ca",	x"06c2",	x"06c4",	x"06fc",	
												x"06e0",	x"06dd",	x"06a1",	x"0706",	
												x"06c8",	x"06fa",	x"06d8",	x"0701",	
												x"06f4",	x"070d",	x"06ed",	x"0708",	
												x"06d8",	x"06f9",	x"06cb",	x"06ee",	
												x"06cb",	x"06c7",	x"06af",	x"06cd",	
												x"06ed",	x"06c1",	x"06d7",	x"06f4",	
												x"06da",	x"06d0",	x"06e1",	x"06d5",	
												x"06db",	x"06ca",	x"06fc",	x"06e1",	
												x"06ff",	x"0707",	x"069c",	x"06f3",	
												x"06c0",	x"06bb",	x"06db",	x"06d2",	
												x"06e3",	x"06d0",	x"06e9",	x"06e4",	
												x"06f1",	x"06e7",	x"0724",	x"06f0",	
												x"0703",	x"0706",	x"068b",	x"06ef",	
												x"3030",	x"3257",	x"0684",	x"06a5",	
												x"0690",	x"0695",	x"0698",	x"0697",	
												x"069d",	x"069a",	x"06be",	x"0692",	
												x"06cb",	x"0688",	x"06bc",	x"06dc",	
												x"06a2",	x"06cf",	x"06da",	x"06e4",	
												x"06c0",	x"06c8",	x"06ce",	x"06c8",	
												x"06cc",	x"06c8",	x"06d0",	x"06ce",	
												x"06ad",	x"06ce",	x"06a8",	x"06b7",	
												x"0693",	x"06ac",	x"06af",	x"06bb",	
												x"06d3",	x"06b1",	x"06bf",	x"06b9",	
												x"06c6",	x"06ce",	x"06d8",	x"06c8",	
												x"06e2",	x"06d6",	x"06ea",	x"06e9",	
												x"06b7",	x"06d9",	x"06d0",	x"06b3",	
												x"06d2",	x"06ca",	x"06dc",	x"06d4",	
												x"06fe",	x"06e2",	x"0706",	x"06f0",	
												x"0708",	x"06ea",	x"06f6",	x"06ef",	
												x"06ad",	x"06d5",	x"0004",	x"000a",	
												x"0c06",	x"be9c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"3258",	
												x"06a1",	x"06ad",	x"06b9",	x"069e",	
												x"06a0",	x"068c",	x"069c",	x"06a6",	
												x"06b4",	x"06a3",	x"06c0",	x"06cd",	
												x"06c2",	x"06c7",	x"06bc",	x"06ee",	
												x"06ec",	x"06dd",	x"06e1",	x"06f2",	
												x"06e5",	x"0706",	x"06e9",	x"06ec",	
												x"0709",	x"06ee",	x"06f0",	x"06f5",	
												x"06f6",	x"0701",	x"06c6",	x"06fb",	
												x"06e7",	x"06e3",	x"0700",	x"06f1",	
												x"0701",	x"0724",	x"070c",	x"0734",	
												x"06fe",	x"0706",	x"06f8",	x"06f6",	
												x"070c",	x"0705",	x"06fb",	x"0713",	
												x"071a",	x"071c",	x"0725",	x"0717",	
												x"0728",	x"071d",	x"0734",	x"0727",	
												x"073c",	x"071b",	x"0744",	x"0734",	
												x"0743",	x"0734",	x"06c0",	x"0729",	
												x"5030",	x"3258",	x"06e4",	x"06df",	
												x"06e2",	x"0700",	x"06e0",	x"06aa",	
												x"06f1",	x"06fa",	x"06fb",	x"06f4",	
												x"06f7",	x"0718",	x"0721",	x"0729",	
												x"0718",	x"0730",	x"072e",	x"072d",	
												x"072c",	x"0720",	x"0728",	x"0728",	
												x"0711",	x"0725",	x"0702",	x"071c",	
												x"0718",	x"070f",	x"072e",	x"0714",	
												x"06ff",	x"0713",	x"0730",	x"0717",	
												x"072f",	x"0736",	x"072d",	x"0736",	
												x"0747",	x"0717",	x"0750",	x"0710",	
												x"0769",	x"0736",	x"0758",	x"0749",	
												x"0735",	x"073e",	x"0745",	x"0723",	
												x"073b",	x"073e",	x"0754",	x"073f",	
												x"077a",	x"073e",	x"0784",	x"0750",	
												x"0772",	x"0753",	x"0769",	x"074d",	
												x"0704",	x"0735",	x"6030",	x"3258",	
												x"070b",	x"0702",	x"06f2",	x"06d7",	
												x"06f4",	x"06e5",	x"0728",	x"06d0",	
												x"0725",	x"070e",	x"071d",	x"072c",	
												x"0731",	x"072d",	x"0740",	x"0733",	
												x"0748",	x"0732",	x"0761",	x"072e",	
												x"074b",	x"073d",	x"075a",	x"075a",	
												x"0750",	x"073c",	x"0748",	x"0748",	
												x"076d",	x"074f",	x"0733",	x"074d",	
												x"0758",	x"0747",	x"0763",	x"0757",	
												x"075c",	x"074f",	x"0776",	x"0747",	
												x"0774",	x"0763",	x"0796",	x"0781",	
												x"077c",	x"0767",	x"0753",	x"076d",	
												x"0795",	x"0759",	x"078b",	x"0768",	
												x"07a7",	x"0761",	x"07a1",	x"0782",	
												x"07b0",	x"0778",	x"07ae",	x"0795",	
												x"07ac",	x"0796",	x"0741",	x"0779",	
												x"7030",	x"3258",	x"0736",	x"0755",	
												x"0764",	x"0732",	x"076e",	x"0750",	
												x"0783",	x"076a",	x"0769",	x"074b",	
												x"0798",	x"0739",	x"07a1",	x"0787",	
												x"0782",	x"0797",	x"07cc",	x"0760",	
												x"07dc",	x"07cc",	x"07a4",	x"07d0",	
												x"07cf",	x"07c1",	x"07c4",	x"07b8",	
												x"07e6",	x"07bb",	x"07e9",	x"07c0",	
												x"07a0",	x"07e6",	x"07e0",	x"07b5",	
												x"07df",	x"07bc",	x"07d1",	x"07df",	
												x"07fb",	x"07d4",	x"07ef",	x"07ee",	
												x"07f0",	x"07ea",	x"0807",	x"07ff",	
												x"07e2",	x"0807",	x"0808",	x"07e2",	
												x"0808",	x"0807",	x"0807",	x"07fb",	
												x"083b",	x"0813",	x"0836",	x"0817",	
												x"083c",	x"0818",	x"0817",	x"082b",	
												x"0761",	x"0814",	x"0004",	x"000a",	
												x"47e0",	x"f13e",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"0259",	
												x"079a",	x"0796",	x"0789",	x"078b",	
												x"0767",	x"0778",	x"07a0",	x"0763",	
												x"077c",	x"077e",	x"077c",	x"0780",	
												x"0740",	x"0778",	x"0721",	x"0754",	
												x"0732",	x"0744",	x"0740",	x"0735",	
												x"073f",	x"072b",	x"072f",	x"0758",	
												x"0744",	x"0732",	x"0779",	x"0760",	
												x"073a",	x"0789",	x"075c",	x"0777",	
												x"077d",	x"077b",	x"078e",	x"079a",	
												x"0784",	x"0778",	x"079e",	x"07a1",	
												x"077e",	x"0769",	x"077d",	x"0785",	
												x"076c",	x"0776",	x"074f",	x"076a",	
												x"076e",	x"0760",	x"0773",	x"0772",	
												x"075a",	x"0757",	x"0764",	x"0777",	
												x"0761",	x"076a",	x"0760",	x"0742",	
												x"0767",	x"0766",	x"071a",	x"075d",	
												x"1031",	x"0259",	x"0748",	x"0763",	
												x"0737",	x"0763",	x"0749",	x"0775",	
												x"0763",	x"0762",	x"074f",	x"075e",	
												x"0748",	x"075f",	x"072e",	x"073c",	
												x"070c",	x"0739",	x"070e",	x"0708",	
												x"0720",	x"070d",	x"0709",	x"070e",	
												x"0755",	x"0726",	x"0725",	x"073a",	
												x"0740",	x"0737",	x"0748",	x"0725",	
												x"0759",	x"0753",	x"0744",	x"0740",	
												x"0778",	x"0761",	x"0778",	x"076c",	
												x"0760",	x"0778",	x"0760",	x"0778",	
												x"0778",	x"0779",	x"0751",	x"0775",	
												x"071d",	x"0752",	x"0741",	x"0743",	
												x"0740",	x"0755",	x"0747",	x"0756",	
												x"077d",	x"0755",	x"0791",	x"0777",	
												x"0778",	x"0770",	x"0768",	x"077b",	
												x"072f",	x"0774",	x"2031",	x"0259",	
												x"074b",	x"0744",	x"0744",	x"074c",	
												x"0753",	x"075f",	x"074a",	x"074f",	
												x"072d",	x"0742",	x"070d",	x"0723",	
												x"072d",	x"070f",	x"06f8",	x"0734",	
												x"072d",	x"0723",	x"0709",	x"0720",	
												x"0706",	x"0707",	x"0705",	x"0742",	
												x"0731",	x"072c",	x"0726",	x"0724",	
												x"0736",	x"0740",	x"0732",	x"0754",	
												x"0785",	x"0742",	x"075b",	x"076c",	
												x"0752",	x"0761",	x"0759",	x"075f",	
												x"0750",	x"0732",	x"074d",	x"0739",	
												x"075a",	x"0741",	x"071d",	x"0745",	
												x"0764",	x"073c",	x"0750",	x"0745",	
												x"0742",	x"0760",	x"0743",	x"0745",	
												x"074c",	x"074b",	x"0759",	x"0741",	
												x"0743",	x"0741",	x"0710",	x"0737",	
												x"3031",	x"0259",	x"0722",	x"070b",	
												x"072d",	x"0723",	x"072d",	x"0723",	
												x"071c",	x"0711",	x"0734",	x"0715",	
												x"0728",	x"0722",	x"06f8",	x"0705",	
												x"06f2",	x"06f1",	x"0705",	x"06d9",	
												x"06f8",	x"0720",	x"070e",	x"06d3",	
												x"06ed",	x"0705",	x"0707",	x"0707",	
												x"072c",	x"0727",	x"0725",	x"073c",	
												x"072a",	x"0723",	x"072f",	x"072a",	
												x"0747",	x"073a",	x"074c",	x"0757",	
												x"0754",	x"073d",	x"0739",	x"0751",	
												x"0740",	x"0731",	x"0744",	x"073b",	
												x"0710",	x"0724",	x"0747",	x"0703",	
												x"074e",	x"0741",	x"074e",	x"0729",	
												x"0760",	x"0756",	x"074d",	x"0743",	
												x"0744",	x"072f",	x"075a",	x"073b",	
												x"0715",	x"0735",	x"0004",	x"000a",	
												x"4240",	x"3153",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"025a",	
												x"0742",	x"074e",	x"0739",	x"0735",	
												x"0745",	x"0734",	x"0740",	x"0745",	
												x"0732",	x"0726",	x"0748",	x"072d",	
												x"072f",	x"072c",	x"0703",	x"072e",	
												x"0727",	x"070a",	x"0716",	x"0705",	
												x"072b",	x"070f",	x"0735",	x"071f",	
												x"0761",	x"072a",	x"075c",	x"075f",	
												x"0769",	x"0764",	x"0768",	x"0776",	
												x"0783",	x"0766",	x"078e",	x"078c",	
												x"0787",	x"0780",	x"0782",	x"0777",	
												x"0774",	x"0792",	x"0791",	x"0793",	
												x"0779",	x"0780",	x"076e",	x"076a",	
												x"07ac",	x"0773",	x"079c",	x"0784",	
												x"077b",	x"0783",	x"0791",	x"079d",	
												x"079b",	x"0793",	x"0793",	x"077c",	
												x"0796",	x"0772",	x"076c",	x"076f",	
												x"5031",	x"025a",	x"0789",	x"0776",	
												x"0767",	x"0767",	x"0780",	x"076d",	
												x"0788",	x"076a",	x"0773",	x"0754",	
												x"0768",	x"0767",	x"0782",	x"075c",	
												x"0757",	x"0754",	x"0767",	x"0762",	
												x"076b",	x"0755",	x"0770",	x"0764",	
												x"077e",	x"0779",	x"0794",	x"0778",	
												x"079b",	x"078e",	x"079c",	x"0781",	
												x"07a2",	x"078a",	x"07b5",	x"0787",	
												x"07c5",	x"0796",	x"079f",	x"0768",	
												x"07ca",	x"0798",	x"07d3",	x"07bd",	
												x"07c6",	x"07ab",	x"07c4",	x"079a",	
												x"07bc",	x"07a7",	x"07d7",	x"077d",	
												x"07c8",	x"078f",	x"07d3",	x"0792",	
												x"07d6",	x"0784",	x"07ea",	x"078c",	
												x"07ec",	x"07ab",	x"07e6",	x"07b7",	
												x"077f",	x"07ac",	x"6031",	x"025a",	
												x"079b",	x"0775",	x"079e",	x"0778",	
												x"079a",	x"0791",	x"0799",	x"0777",	
												x"079f",	x"0779",	x"07a2",	x"0782",	
												x"078b",	x"0781",	x"075f",	x"0750",	
												x"0783",	x"0746",	x"0788",	x"0773",	
												x"0794",	x"075d",	x"07b2",	x"078e",	
												x"07c5",	x"077d",	x"07d5",	x"07ad",	
												x"07df",	x"07b2",	x"07cb",	x"07bd",	
												x"0805",	x"07bc",	x"07f3",	x"07f2",	
												x"07f6",	x"07e0",	x"0816",	x"07ee",	
												x"07fa",	x"07e5",	x"07f7",	x"07d4",	
												x"081e",	x"07e7",	x"07e3",	x"07f2",	
												x"081c",	x"07b5",	x"0815",	x"0803",	
												x"07f7",	x"07da",	x"0807",	x"07d2",	
												x"081f",	x"07de",	x"0823",	x"0800",	
												x"0816",	x"07e6",	x"07ee",	x"07d6",	
												x"7031",	x"025a",	x"07fc",	x"07f8",	
												x"0811",	x"07cd",	x"0809",	x"07d5",	
												x"081d",	x"07e6",	x"0814",	x"0800",	
												x"0821",	x"07f4",	x"07fe",	x"07b3",	
												x"07e2",	x"07bd",	x"07c5",	x"07b2",	
												x"07d3",	x"07d6",	x"07ea",	x"07c5",	
												x"083a",	x"07e6",	x"080c",	x"07ce",	
												x"082c",	x"07ef",	x"084c",	x"0823",	
												x"0861",	x"0842",	x"0868",	x"081b",	
												x"0866",	x"0854",	x"0875",	x"0850",	
												x"088e",	x"085e",	x"085b",	x"0876",	
												x"088d",	x"0867",	x"087c",	x"0883",	
												x"087c",	x"0878",	x"0884",	x"0878",	
												x"089d",	x"0875",	x"089b",	x"087f",	
												x"08d4",	x"089b",	x"08b4",	x"086a",	
												x"08be",	x"088e",	x"089c",	x"089e",	
												x"05f8",	x"089c",	x"0004",	x"000a",	
												x"8220",	x"6457",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"125b",	
												x"05e7",	x"05fc",	x"05fd",	x"05fb",	
												x"05c0",	x"05f7",	x"05d5",	x"05d7",	
												x"05b9",	x"05d3",	x"05e6",	x"05df",	
												x"05aa",	x"05db",	x"05c8",	x"05cd",	
												x"05df",	x"05e2",	x"0604",	x"05f5",	
												x"05fe",	x"05ff",	x"0627",	x"060e",	
												x"0619",	x"0636",	x"0614",	x"0633",	
												x"061b",	x"0641",	x"060b",	x"0616",	
												x"0612",	x"0607",	x"060d",	x"062b",	
												x"0604",	x"0611",	x"0605",	x"0610",	
												x"0601",	x"0612",	x"0624",	x"0605",	
												x"060c",	x"0603",	x"060a",	x"0616",	
												x"0600",	x"05fc",	x"0620",	x"060d",	
												x"0613",	x"061d",	x"0613",	x"0634",	
												x"063b",	x"0607",	x"0644",	x"0629",	
												x"062a",	x"0622",	x"05df",	x"0616",	
												x"1031",	x"125b",	x"05e8",	x"05eb",	
												x"05dc",	x"05e7",	x"05ea",	x"05df",	
												x"05be",	x"05dd",	x"05ca",	x"05ab",	
												x"05a0",	x"05b0",	x"05d4",	x"05a7",	
												x"05be",	x"05e9",	x"05e1",	x"05cf",	
												x"0607",	x"05fb",	x"0614",	x"05f2",	
												x"0631",	x"0608",	x"05fe",	x"0613",	
												x"05fa",	x"05fe",	x"05f9",	x"060d",	
												x"05cf",	x"0615",	x"05f3",	x"05ee",	
												x"0603",	x"05fd",	x"0609",	x"0616",	
												x"05fd",	x"0611",	x"05fd",	x"060a",	
												x"0601",	x"060d",	x"05f7",	x"060a",	
												x"05d1",	x"0610",	x"060d",	x"05f8",	
												x"0603",	x"05fb",	x"0617",	x"0621",	
												x"0604",	x"061c",	x"061c",	x"060c",	
												x"0622",	x"0620",	x"0614",	x"061f",	
												x"05b8",	x"060b",	x"2031",	x"125b",	
												x"05cd",	x"05ea",	x"05e0",	x"05e4",	
												x"05c0",	x"05cc",	x"05c9",	x"05c8",	
												x"05b6",	x"05ae",	x"05ab",	x"05d3",	
												x"05c7",	x"05d1",	x"05bb",	x"05dd",	
												x"05c1",	x"05d0",	x"05e7",	x"05db",	
												x"05fc",	x"05f0",	x"05ec",	x"05e4",	
												x"0616",	x"05ef",	x"05f2",	x"060b",	
												x"05ec",	x"05ef",	x"05dd",	x"05fe",	
												x"05e6",	x"05dc",	x"05e3",	x"05ea",	
												x"0606",	x"05fa",	x"0600",	x"0609",	
												x"0603",	x"05e8",	x"05ff",	x"0601",	
												x"05fc",	x"0601",	x"05be",	x"0600",	
												x"05f4",	x"05e6",	x"05fb",	x"05f8",	
												x"0603",	x"05e8",	x"0614",	x"0607",	
												x"0611",	x"0603",	x"0607",	x"0611",	
												x"0613",	x"0601",	x"05d3",	x"05f6",	
												x"3031",	x"125b",	x"05a8",	x"05be",	
												x"05ad",	x"05ae",	x"05de",	x"05a7",	
												x"05d6",	x"05d4",	x"05c0",	x"05ba",	
												x"05b9",	x"05a1",	x"05c2",	x"05aa",	
												x"05ac",	x"059c",	x"05e5",	x"05c2",	
												x"05e8",	x"05dc",	x"05f5",	x"05dd",	
												x"05fd",	x"05fa",	x"05fa",	x"05f2",	
												x"0600",	x"05f1",	x"05f8",	x"05f1",	
												x"05cb",	x"05f3",	x"0609",	x"05b3",	
												x"0610",	x"05f3",	x"060e",	x"05f8",	
												x"0615",	x"05f8",	x"060d",	x"060f",	
												x"060d",	x"0602",	x"0621",	x"05f6",	
												x"05eb",	x"05e7",	x"0624",	x"05e3",	
												x"0615",	x"05fc",	x"0627",	x"05f4",	
												x"0623",	x"0614",	x"0627",	x"05ff",	
												x"0631",	x"060f",	x"062f",	x"0611",	
												x"05de",	x"05ff",	x"0004",	x"000a",	
												x"99c1",	x"c76a",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"125c",	
												x"05f7",	x"05d6",	x"05fe",	x"05db",	
												x"05e9",	x"05e7",	x"05e5",	x"05d4",	
												x"05e3",	x"05c7",	x"05e5",	x"05cd",	
												x"05d8",	x"05cf",	x"05ee",	x"05d5",	
												x"05f2",	x"05c9",	x"060d",	x"05eb",	
												x"0637",	x"0614",	x"0621",	x"0627",	
												x"0626",	x"0614",	x"062e",	x"062b",	
												x"0639",	x"0610",	x"0606",	x"061e",	
												x"0638",	x"0619",	x"063a",	x"062d",	
												x"0645",	x"0635",	x"0650",	x"0639",	
												x"0649",	x"063e",	x"063f",	x"063a",	
												x"0633",	x"0632",	x"062d",	x"0632",	
												x"0652",	x"0627",	x"0659",	x"0645",	
												x"064b",	x"0639",	x"0650",	x"0644",	
												x"065a",	x"0644",	x"0659",	x"0653",	
												x"0662",	x"0658",	x"0616",	x"0641",	
												x"5031",	x"125c",	x"0640",	x"05fe",	
												x"0625",	x"0618",	x"0624",	x"05d7",	
												x"060b",	x"0602",	x"0623",	x"0609",	
												x"0629",	x"0615",	x"0630",	x"060a",	
												x"061f",	x"0603",	x"065d",	x"061d",	
												x"0666",	x"0646",	x"0648",	x"0648",	
												x"0658",	x"064c",	x"065f",	x"063a",	
												x"0655",	x"065a",	x"0654",	x"061f",	
												x"0650",	x"0638",	x"0669",	x"063a",	
												x"0673",	x"0652",	x"0673",	x"063b",	
												x"0671",	x"064e",	x"068f",	x"0651",	
												x"0691",	x"065a",	x"0678",	x"064e",	
												x"0671",	x"0657",	x"0680",	x"0657",	
												x"069b",	x"065d",	x"0683",	x"0648",	
												x"06b4",	x"065e",	x"06ac",	x"0659",	
												x"0699",	x"066d",	x"0683",	x"0678",	
												x"0633",	x"0668",	x"6031",	x"125c",	
												x"062e",	x"062a",	x"0642",	x"0616",	
												x"0636",	x"0618",	x"0642",	x"0623",	
												x"0647",	x"0625",	x"0634",	x"0626",	
												x"0641",	x"061f",	x"063d",	x"060f",	
												x"0663",	x"0615",	x"0666",	x"061d",	
												x"0681",	x"0651",	x"0685",	x"0662",	
												x"068f",	x"065e",	x"0697",	x"0670",	
												x"0688",	x"067d",	x"0673",	x"0688",	
												x"0690",	x"0661",	x"0681",	x"068f",	
												x"06a1",	x"066e",	x"06a4",	x"0687",	
												x"06b6",	x"0693",	x"06a3",	x"0682",	
												x"06b0",	x"0688",	x"068d",	x"0691",	
												x"06ab",	x"067a",	x"06b6",	x"067b",	
												x"06cf",	x"0693",	x"06c6",	x"0699",	
												x"06c8",	x"068b",	x"06c8",	x"069d",	
												x"06b4",	x"0697",	x"0691",	x"067e",	
												x"7031",	x"125c",	x"068b",	x"0659",	
												x"0687",	x"0659",	x"0675",	x"062d",	
												x"069e",	x"0648",	x"0697",	x"064b",	
												x"068c",	x"0640",	x"06a6",	x"0661",	
												x"0683",	x"0668",	x"06e5",	x"0664",	
												x"06e3",	x"068f",	x"06e5",	x"06a8",	
												x"06e3",	x"06cf",	x"06f3",	x"069a",	
												x"06f0",	x"06e8",	x"06ee",	x"06e1",	
												x"06c1",	x"06c1",	x"070b",	x"06c1",	
												x"071a",	x"06d5",	x"070d",	x"06de",	
												x"0700",	x"06e3",	x"0721",	x"06ef",	
												x"0720",	x"0701",	x"0714",	x"06fe",	
												x"06f9",	x"06ed",	x"071b",	x"06f1",	
												x"0729",	x"0714",	x"0724",	x"0709",	
												x"0739",	x"071d",	x"0754",	x"0718",	
												x"073e",	x"070e",	x"073c",	x"071b",	
												x"06c8",	x"0712",	x"0004",	x"000a",	
												x"de0d",	x"fb3f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"225d",	
												x"06e2",	x"0705",	x"06c8",	x"06c4",	
												x"06b2",	x"06a8",	x"06b5",	x"06b2",	
												x"06c1",	x"06ac",	x"06ed",	x"06de",	
												x"06d1",	x"06e9",	x"06b8",	x"06db",	
												x"06dc",	x"06c5",	x"06e4",	x"06ff",	
												x"06ea",	x"06fd",	x"070b",	x"071e",	
												x"06f4",	x"0709",	x"0716",	x"0721",	
												x"06d9",	x"0725",	x"06df",	x"06ed",	
												x"06de",	x"0706",	x"06f2",	x"06f2",	
												x"06f5",	x"06ed",	x"0712",	x"06fc",	
												x"06f3",	x"070a",	x"06eb",	x"0707",	
												x"06d8",	x"0700",	x"06e3",	x"06f5",	
												x"071f",	x"06f0",	x"06f2",	x"0712",	
												x"06ea",	x"06dc",	x"072c",	x"06fe",	
												x"070b",	x"06ef",	x"0730",	x"0708",	
												x"06e1",	x"06d5",	x"0696",	x"06c9",	
												x"1031",	x"225d",	x"06b5",	x"06bc",	
												x"06dd",	x"06d1",	x"06b8",	x"06d6",	
												x"069a",	x"06bb",	x"06d3",	x"06a1",	
												x"06be",	x"06bf",	x"06c5",	x"0692",	
												x"06c4",	x"06c6",	x"06d0",	x"06ce",	
												x"070d",	x"06f6",	x"06f4",	x"06f6",	
												x"06ee",	x"06ed",	x"06e6",	x"06ec",	
												x"06ca",	x"06ee",	x"06d3",	x"06eb",	
												x"0696",	x"06ca",	x"06cf",	x"06ce",	
												x"06e6",	x"06d7",	x"06e4",	x"06f8",	
												x"06e2",	x"06ed",	x"06f3",	x"06e4",	
												x"06e4",	x"06eb",	x"06cd",	x"06e7",	
												x"06b0",	x"06e8",	x"06d7",	x"06ef",	
												x"070a",	x"06e8",	x"06e5",	x"0712",	
												x"0717",	x"06fd",	x"070d",	x"06f0",	
												x"06fe",	x"0704",	x"06ea",	x"0701",	
												x"0691",	x"070e",	x"2031",	x"225d",	
												x"06b0",	x"06c8",	x"06bb",	x"06a7",	
												x"06a3",	x"06d3",	x"06a0",	x"06be",	
												x"067d",	x"0696",	x"068f",	x"0686",	
												x"0693",	x"0698",	x"0689",	x"06ad",	
												x"06d2",	x"06b4",	x"06cd",	x"06e7",	
												x"06df",	x"06f1",	x"06b6",	x"06d3",	
												x"06cf",	x"06c7",	x"06db",	x"06fe",	
												x"06d0",	x"06d5",	x"06c8",	x"06d7",	
												x"06ce",	x"06d4",	x"06d5",	x"06cb",	
												x"06e5",	x"06e2",	x"06db",	x"06e1",	
												x"06f8",	x"06e3",	x"06e0",	x"06e7",	
												x"06e3",	x"06d4",	x"06bb",	x"06ec",	
												x"06e0",	x"06ac",	x"06d8",	x"06dc",	
												x"06ec",	x"06d7",	x"06ed",	x"06f4",	
												x"06fb",	x"06da",	x"06fa",	x"06e5",	
												x"06f3",	x"06eb",	x"0694",	x"06e5",	
												x"3031",	x"225d",	x"06b6",	x"068a",	
												x"06a1",	x"066c",	x"0681",	x"0669",	
												x"0690",	x"0684",	x"06c8",	x"066b",	
												x"06a1",	x"068e",	x"06ab",	x"0697",	
												x"0680",	x"06ae",	x"068e",	x"0687",	
												x"06d2",	x"06b0",	x"06ab",	x"06d4",	
												x"06b3",	x"06af",	x"06e1",	x"06b6",	
												x"06dc",	x"06ba",	x"06c4",	x"06c9",	
												x"06ae",	x"06c7",	x"06a7",	x"06b2",	
												x"06df",	x"06b9",	x"06ef",	x"06c8",	
												x"070e",	x"06e0",	x"06e3",	x"06c7",	
												x"06d0",	x"06cf",	x"06dc",	x"06c3",	
												x"06e5",	x"06c7",	x"06f2",	x"06c4",	
												x"06dd",	x"06c0",	x"06e9",	x"06db",	
												x"0705",	x"06d4",	x"0712",	x"06dd",	
												x"0711",	x"06db",	x"06fb",	x"06e9",	
												x"06d5",	x"06da",	x"0004",	x"000a",	
												x"0a72",	x"781f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"225e",	
												x"06a7",	x"069b",	x"06a6",	x"0689",	
												x"06a4",	x"0687",	x"06dd",	x"06a0",	
												x"06cd",	x"0692",	x"06c9",	x"06aa",	
												x"06bf",	x"06d8",	x"06a5",	x"06af",	
												x"06fe",	x"06d0",	x"0704",	x"06d7",	
												x"06ee",	x"06e9",	x"06ff",	x"06d0",	
												x"0711",	x"06f3",	x"0714",	x"0707",	
												x"0709",	x"0703",	x"070d",	x"0711",	
												x"0711",	x"06f1",	x"0718",	x"0713",	
												x"0710",	x"071e",	x"071e",	x"06fd",	
												x"0723",	x"070b",	x"072a",	x"0721",	
												x"0724",	x"071d",	x"0718",	x"0701",	
												x"0730",	x"0713",	x"0739",	x"0724",	
												x"073c",	x"0710",	x"0751",	x"0722",	
												x"074e",	x"0731",	x"0750",	x"0730",	
												x"074e",	x"0714",	x"06f6",	x"0717",	
												x"5031",	x"225e",	x"070c",	x"06ce",	
												x"06ff",	x"06f1",	x"06e0",	x"06ea",	
												x"06fb",	x"06d1",	x"0720",	x"06ef",	
												x"0709",	x"06fe",	x"0724",	x"06fa",	
												x"0700",	x"0710",	x"0720",	x"06d9",	
												x"0746",	x"06fc",	x"0741",	x"0729",	
												x"072d",	x"071c",	x"073d",	x"0729",	
												x"0744",	x"0729",	x"0752",	x"071e",	
												x"0730",	x"0719",	x"0747",	x"071d",	
												x"0756",	x"0727",	x"074f",	x"073e",	
												x"0746",	x"0733",	x"0760",	x"072e",	
												x"075b",	x"0733",	x"0756",	x"072c",	
												x"075d",	x"073a",	x"0772",	x"06f8",	
												x"077b",	x"0738",	x"0770",	x"0735",	
												x"0772",	x"0740",	x"077d",	x"0745",	
												x"0768",	x"0737",	x"0771",	x"0740",	
												x"06f5",	x"0741",	x"6031",	x"225e",	
												x"074d",	x"06eb",	x"06f8",	x"06dd",	
												x"070b",	x"06d2",	x"0723",	x"06dd",	
												x"071c",	x"0706",	x"0728",	x"06fa",	
												x"072d",	x"0706",	x"0745",	x"071c",	
												x"0757",	x"0713",	x"076d",	x"0745",	
												x"075c",	x"0753",	x"076e",	x"0753",	
												x"078e",	x"0727",	x"07a2",	x"0762",	
												x"0794",	x"0757",	x"0767",	x"0764",	
												x"0782",	x"074f",	x"0783",	x"078a",	
												x"0795",	x"075e",	x"0795",	x"075c",	
												x"0796",	x"076b",	x"07a0",	x"075e",	
												x"0791",	x"0773",	x"0785",	x"0759",	
												x"07a0",	x"0769",	x"07b1",	x"0764",	
												x"07cb",	x"076b",	x"07c1",	x"0785",	
												x"07c3",	x"0787",	x"07b8",	x"0776",	
												x"07a7",	x"0783",	x"0733",	x"078c",	
												x"7031",	x"225e",	x"075d",	x"073d",	
												x"0765",	x"0748",	x"0736",	x"0740",	
												x"0797",	x"0733",	x"0781",	x"0741",	
												x"075b",	x"072f",	x"0761",	x"0748",	
												x"078e",	x"0761",	x"07cd",	x"077c",	
												x"07bb",	x"0798",	x"07ec",	x"07be",	
												x"07f5",	x"07c8",	x"0803",	x"07d4",	
												x"07ff",	x"07d3",	x"07df",	x"07b2",	
												x"07ad",	x"07c0",	x"0812",	x"07ae",	
												x"0831",	x"07e9",	x"07fb",	x"07e3",	
												x"0841",	x"07fd",	x"081f",	x"07dc",	
												x"0809",	x"07ec",	x"0829",	x"0801",	
												x"07e9",	x"07e4",	x"0834",	x"07d3",	
												x"0825",	x"0819",	x"0824",	x"081b",	
												x"083e",	x"081e",	x"085e",	x"081a",	
												x"084b",	x"0833",	x"0835",	x"0831",	
												x"06da",	x"0828",	x"0004",	x"000a",	
												x"521a",	x"aef3",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"325f",	
												x"06b8",	x"06e0",	x"06c0",	x"06b8",	
												x"06b8",	x"06c0",	x"06b4",	x"06bc",	
												x"06b1",	x"06b3",	x"06cd",	x"06b1",	
												x"0709",	x"06ca",	x"06cc",	x"06d2",	
												x"06e4",	x"06eb",	x"070d",	x"06eb",	
												x"06fa",	x"06fd",	x"0720",	x"06fa",	
												x"06f5",	x"071d",	x"070b",	x"0719",	
												x"072d",	x"071f",	x"06a2",	x"0718",	
												x"06da",	x"06d5",	x"0709",	x"06f1",	
												x"0710",	x"0710",	x"0704",	x"0721",	
												x"0715",	x"06f6",	x"06fe",	x"0728",	
												x"06ef",	x"070d",	x"06fe",	x"071d",	
												x"0730",	x"06fc",	x"072e",	x"0738",	
												x"071c",	x"0700",	x"0702",	x"0711",	
												x"06ef",	x"06ee",	x"0726",	x"06f9",	
												x"0703",	x"070b",	x"06ab",	x"06f7",	
												x"1031",	x"325f",	x"06b0",	x"06b9",	
												x"06bb",	x"06c1",	x"06ae",	x"06d2",	
												x"06ab",	x"06f1",	x"06aa",	x"06a3",	
												x"06b3",	x"06a8",	x"06c2",	x"06d7",	
												x"06a1",	x"06d6",	x"06eb",	x"06eb",	
												x"06e2",	x"06eb",	x"06e7",	x"06f0",	
												x"06f8",	x"06f5",	x"06e6",	x"06ef",	
												x"06e5",	x"070b",	x"070e",	x"06e7",	
												x"069f",	x"06eb",	x"06bf",	x"06d1",	
												x"06ed",	x"06e3",	x"06ec",	x"06e5",	
												x"06e4",	x"070d",	x"06e4",	x"06e5",	
												x"0702",	x"0703",	x"06e6",	x"0716",	
												x"06b6",	x"06f1",	x"0702",	x"0711",	
												x"071d",	x"06eb",	x"071c",	x"0700",	
												x"06f8",	x"06f6",	x"0702",	x"06eb",	
												x"0707",	x"06ee",	x"070d",	x"0714",	
												x"06b5",	x"070c",	x"2031",	x"325f",	
												x"06a7",	x"06c2",	x"06a5",	x"06a0",	
												x"06ae",	x"0699",	x"069f",	x"06bd",	
												x"06b6",	x"06cd",	x"06c7",	x"06d9",	
												x"06e0",	x"06d0",	x"069d",	x"06e9",	
												x"06d5",	x"06d2",	x"06e4",	x"06f5",	
												x"06cd",	x"0708",	x"06c3",	x"06e6",	
												x"06d7",	x"06da",	x"06bf",	x"06ed",	
												x"06ea",	x"06db",	x"06b0",	x"06ea",	
												x"06d9",	x"06b6",	x"06f5",	x"06cb",	
												x"06f6",	x"06d4",	x"06df",	x"06e6",	
												x"06eb",	x"06bb",	x"06ec",	x"06fb",	
												x"06ed",	x"06e3",	x"06e0",	x"06da",	
												x"06ed",	x"06e2",	x"06e9",	x"06e3",	
												x"06eb",	x"06d6",	x"06f3",	x"0706",	
												x"06eb",	x"06cb",	x"06f8",	x"06b8",	
												x"070c",	x"06e7",	x"0681",	x"06d2",	
												x"3031",	x"325f",	x"069a",	x"068e",	
												x"06b2",	x"06ab",	x"0683",	x"068e",	
												x"068e",	x"0682",	x"06c0",	x"0684",	
												x"06c0",	x"0699",	x"06ad",	x"06ac",	
												x"0682",	x"06b6",	x"06e2",	x"06b5",	
												x"06ba",	x"06ce",	x"06c7",	x"06c2",	
												x"06cf",	x"06cc",	x"06da",	x"06da",	
												x"06e1",	x"06d9",	x"06d9",	x"06dc",	
												x"06b5",	x"06dd",	x"06cf",	x"06c5",	
												x"06e2",	x"06ba",	x"06e0",	x"06c9",	
												x"06f0",	x"06fe",	x"06e9",	x"06fe",	
												x"06f9",	x"06e6",	x"06e7",	x"06eb",	
												x"06e2",	x"06e4",	x"06fd",	x"06d8",	
												x"06ed",	x"06e7",	x"06f2",	x"06e8",	
												x"0715",	x"06f1",	x"0719",	x"06f1",	
												x"0718",	x"06ee",	x"06fb",	x"06e0",	
												x"06d5",	x"06db",	x"0004",	x"000a",	
												x"0ea7",	x"bdb5",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"3260",	
												x"06c5",	x"06b5",	x"06a7",	x"06a9",	
												x"06c1",	x"06b2",	x"06a9",	x"06b2",	
												x"06c3",	x"06af",	x"06c6",	x"06d0",	
												x"06cf",	x"06c4",	x"06a4",	x"06e0",	
												x"06f3",	x"06c6",	x"06fd",	x"06df",	
												x"070d",	x"070a",	x"070c",	x"070c",	
												x"070e",	x"06e2",	x"070d",	x"06ea",	
												x"0703",	x"06f5",	x"06fd",	x"0701",	
												x"0718",	x"06ff",	x"0729",	x"0714",	
												x"072d",	x"073f",	x"073a",	x"0714",	
												x"0739",	x"0721",	x"0739",	x"0724",	
												x"0737",	x"0723",	x"0714",	x"071b",	
												x"0739",	x"0723",	x"073d",	x"072a",	
												x"072f",	x"072a",	x"0724",	x"072f",	
												x"0726",	x"0705",	x"0759",	x"0716",	
												x"0760",	x"0723",	x"06f4",	x"0720",	
												x"5031",	x"3260",	x"0701",	x"06fb",	
												x"0708",	x"06e5",	x"0703",	x"06d7",	
												x"0739",	x"06f5",	x"0718",	x"06ec",	
												x"0717",	x"0702",	x"072c",	x"06fe",	
												x"0721",	x"0712",	x"073c",	x"0720",	
												x"0743",	x"072b",	x"0751",	x"0745",	
												x"0748",	x"0743",	x"0756",	x"0739",	
												x"074d",	x"0725",	x"0740",	x"0738",	
												x"0727",	x"072d",	x"0737",	x"071d",	
												x"0755",	x"0740",	x"075a",	x"071f",	
												x"0766",	x"0735",	x"077e",	x"0716",	
												x"0783",	x"074e",	x"0781",	x"0740",	
												x"0762",	x"0738",	x"0796",	x"0732",	
												x"0771",	x"0757",	x"0768",	x"0743",	
												x"077a",	x"0741",	x"0799",	x"0752",	
												x"0795",	x"0759",	x"077c",	x"075a",	
												x"06ea",	x"074c",	x"6031",	x"3260",	
												x"0736",	x"06ed",	x"0713",	x"06f0",	
												x"0729",	x"06d6",	x"0731",	x"0703",	
												x"073f",	x"06e2",	x"0733",	x"0720",	
												x"073b",	x"071a",	x"0732",	x"0731",	
												x"075a",	x"0715",	x"076f",	x"0729",	
												x"0799",	x"0761",	x"0797",	x"076c",	
												x"076c",	x"074c",	x"0777",	x"0759",	
												x"0784",	x"075c",	x"076c",	x"0767",	
												x"0783",	x"076d",	x"0799",	x"0779",	
												x"079a",	x"077d",	x"07b0",	x"076d",	
												x"07a2",	x"0777",	x"07be",	x"078f",	
												x"07ac",	x"077d",	x"078c",	x"077a",	
												x"079c",	x"0792",	x"07dc",	x"0799",	
												x"07bc",	x"0795",	x"07ac",	x"0791",	
												x"07bb",	x"077e",	x"07d1",	x"0781",	
												x"07d6",	x"0792",	x"075d",	x"0799",	
												x"7031",	x"3260",	x"0783",	x"0729",	
												x"07a0",	x"0744",	x"0771",	x"072a",	
												x"0780",	x"0740",	x"079b",	x"075f",	
												x"079a",	x"077d",	x"07a2",	x"0759",	
												x"077d",	x"075c",	x"07cc",	x"0776",	
												x"07c3",	x"078e",	x"07b5",	x"07b7",	
												x"07cb",	x"07c3",	x"07e2",	x"07bf",	
												x"0814",	x"07dc",	x"0806",	x"07d7",	
												x"07d1",	x"07f6",	x"07ef",	x"07af",	
												x"07fe",	x"07d4",	x"0809",	x"07f2",	
												x"081f",	x"07e1",	x"0819",	x"07f7",	
												x"081a",	x"07f3",	x"082b",	x"07f0",	
												x"081b",	x"07fa",	x"084c",	x"07e8",	
												x"0822",	x"080b",	x"0823",	x"0817",	
												x"0862",	x"0825",	x"085a",	x"0821",	
												x"0870",	x"0821",	x"0836",	x"0835",	
												x"0749",	x"081f",	x"0004",	x"000a",	
												x"5720",	x"f4e5",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"0361",	
												x"0763",	x"0761",	x"074d",	x"0774",	
												x"0741",	x"077a",	x"0748",	x"0740",	
												x"077c",	x"074c",	x"0747",	x"075d",	
												x"0779",	x"0757",	x"076d",	x"075a",	
												x"0797",	x"07a6",	x"0796",	x"07b2",	
												x"07a0",	x"07a6",	x"07b7",	x"07b8",	
												x"0795",	x"07ab",	x"0794",	x"07b6",	
												x"07bc",	x"07b6",	x"078b",	x"0793",	
												x"0777",	x"07a6",	x"07a3",	x"0798",	
												x"07a4",	x"07b2",	x"07ab",	x"07a6",	
												x"0798",	x"07a1",	x"0796",	x"07c2",	
												x"07b6",	x"07bb",	x"072c",	x"0782",	
												x"076c",	x"077d",	x"07c4",	x"07a5",	
												x"07a3",	x"079f",	x"07aa",	x"07ac",	
												x"07a7",	x"07a3",	x"079e",	x"07a4",	
												x"0792",	x"07a9",	x"076c",	x"0765",	
												x"102e",	x"0361",	x"074d",	x"076c",	
												x"0742",	x"075e",	x"0744",	x"0756",	
												x"0740",	x"074e",	x"0742",	x"073c",	
												x"0778",	x"0753",	x"073f",	x"075a",	
												x"0750",	x"0762",	x"0769",	x"076f",	
												x"0785",	x"0775",	x"0794",	x"0784",	
												x"0794",	x"0794",	x"0780",	x"07a6",	
												x"0797",	x"079e",	x"0789",	x"079a",	
												x"0748",	x"0759",	x"0756",	x"076c",	
												x"076f",	x"0787",	x"0795",	x"0784",	
												x"0797",	x"079a",	x"0787",	x"07a9",	
												x"07a4",	x"0790",	x"0768",	x"07a2",	
												x"0750",	x"077e",	x"078b",	x"077e",	
												x"0788",	x"0794",	x"0794",	x"0776",	
												x"07a1",	x"07a5",	x"0797",	x"07b0",	
												x"0787",	x"0790",	x"0799",	x"079b",	
												x"0740",	x"0787",	x"202e",	x"0361",	
												x"0746",	x"0748",	x"073a",	x"0747",	
												x"071f",	x"074a",	x"0724",	x"072a",	
												x"0730",	x"0747",	x"076d",	x"0751",	
												x"0778",	x"076b",	x"0722",	x"0791",	
												x"0765",	x"0761",	x"0760",	x"0783",	
												x"0770",	x"075b",	x"078a",	x"078e",	
												x"075f",	x"0773",	x"0757",	x"0783",	
												x"077d",	x"0772",	x"072c",	x"0776",	
												x"076e",	x"076a",	x"0762",	x"076a",	
												x"0775",	x"0768",	x"0772",	x"0785",	
												x"0777",	x"0773",	x"077f",	x"0780",	
												x"075f",	x"0769",	x"073d",	x"0770",	
												x"0775",	x"077c",	x"078c",	x"0770",	
												x"0774",	x"078b",	x"078f",	x"0791",	
												x"078a",	x"077e",	x"0786",	x"0782",	
												x"0785",	x"0764",	x"070c",	x"0787",	
												x"302e",	x"0361",	x"0715",	x"070a",	
												x"0717",	x"06ef",	x"071f",	x"0721",	
												x"0740",	x"0733",	x"0730",	x"071d",	
												x"072e",	x"0721",	x"0745",	x"0739",	
												x"073d",	x"0755",	x"0730",	x"073b",	
												x"0743",	x"074b",	x"0766",	x"073e",	
												x"0749",	x"0753",	x"0773",	x"0742",	
												x"077b",	x"0778",	x"0754",	x"0747",	
												x"0728",	x"0744",	x"072c",	x"0745",	
												x"074a",	x"074b",	x"075b",	x"0755",	
												x"0774",	x"0755",	x"0772",	x"077f",	
												x"0766",	x"0754",	x"0752",	x"075a",	
												x"073f",	x"0751",	x"0781",	x"0764",	
												x"076b",	x"0763",	x"07ae",	x"075f",	
												x"07b1",	x"079a",	x"0789",	x"0785",	
												x"0792",	x"0777",	x"0791",	x"0765",	
												x"0736",	x"0771",	x"0004",	x"000a",	
												x"55e8",	x"4b1a",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"0362",	
												x"073f",	x"072d",	x"0734",	x"0748",	
												x"0722",	x"0721",	x"0727",	x"070c",	
												x"074f",	x"0722",	x"076d",	x"0755",	
												x"0759",	x"0763",	x"072c",	x"074b",	
												x"0775",	x"0732",	x"0786",	x"076e",	
												x"0782",	x"078e",	x"0787",	x"0788",	
												x"0787",	x"0782",	x"0785",	x"07a3",	
												x"0780",	x"0791",	x"074d",	x"0781",	
												x"079b",	x"076f",	x"07b7",	x"07a0",	
												x"07b5",	x"07a0",	x"07c0",	x"07ae",	
												x"07bc",	x"07b9",	x"07a7",	x"07b7",	
												x"079d",	x"0798",	x"077a",	x"0799",	
												x"07ac",	x"0794",	x"07d0",	x"07b0",	
												x"07d4",	x"07bf",	x"07db",	x"07d6",	
												x"07da",	x"07b9",	x"07d2",	x"07b5",	
												x"07ce",	x"07a4",	x"0797",	x"07aa",	
												x"502e",	x"0362",	x"0784",	x"0760",	
												x"07a2",	x"077c",	x"0765",	x"0762",	
												x"078e",	x"075f",	x"0780",	x"0793",	
												x"0785",	x"0782",	x"0784",	x"0787",	
												x"078d",	x"07ad",	x"07a7",	x"0788",	
												x"07b2",	x"07c2",	x"07d8",	x"07ab",	
												x"07cc",	x"07e1",	x"07e3",	x"07ba",	
												x"07bb",	x"07e2",	x"07c5",	x"07a8",	
												x"0787",	x"079e",	x"07cf",	x"079f",	
												x"07bf",	x"07f0",	x"07d6",	x"079c",	
												x"07f9",	x"07cc",	x"07f0",	x"07e3",	
												x"07e7",	x"07e1",	x"07db",	x"07a9",	
												x"07d2",	x"07d4",	x"07ef",	x"07b5",	
												x"07fe",	x"07bd",	x"0808",	x"07bb",	
												x"0813",	x"07ee",	x"07ff",	x"07ed",	
												x"0808",	x"07ec",	x"07eb",	x"07d9",	
												x"07c1",	x"07da",	x"602e",	x"0362",	
												x"07a2",	x"0784",	x"07b7",	x"079e",	
												x"0792",	x"0782",	x"07b9",	x"0783",	
												x"07c7",	x"0782",	x"07c7",	x"07ba",	
												x"07b1",	x"07a9",	x"07ae",	x"0795",	
												x"07f6",	x"078e",	x"07fc",	x"07d2",	
												x"07ed",	x"07cf",	x"07fd",	x"07eb",	
												x"07f5",	x"07ec",	x"07eb",	x"0816",	
												x"07e7",	x"07e5",	x"07c2",	x"07be",	
												x"07fa",	x"07c2",	x"07f9",	x"0802",	
												x"0806",	x"07f0",	x"0831",	x"07fb",	
												x"081a",	x"0802",	x"0810",	x"07fa",	
												x"0828",	x"07fd",	x"0808",	x"07d1",	
												x"0831",	x"0807",	x"082f",	x"0822",	
												x"084d",	x"081b",	x"0846",	x"0839",	
												x"084f",	x"082e",	x"083d",	x"082a",	
												x"0845",	x"0822",	x"07be",	x"080a",	
												x"702e",	x"0362",	x"07c3",	x"079a",	
												x"07d9",	x"07a9",	x"07b2",	x"07ac",	
												x"07c8",	x"0795",	x"07cf",	x"07cf",	
												x"082e",	x"07c5",	x"07ff",	x"0800",	
												x"07f9",	x"0832",	x"082a",	x"07fc",	
												x"0820",	x"0811",	x"0856",	x"081e",	
												x"086c",	x"085f",	x"0878",	x"086b",	
												x"0860",	x"085c",	x"0846",	x"0855",	
												x"083b",	x"0849",	x"0874",	x"083b",	
												x"087c",	x"0867",	x"087b",	x"086d",	
												x"089e",	x"085c",	x"08ae",	x"0890",	
												x"0896",	x"0890",	x"085a",	x"087e",	
												x"0860",	x"0878",	x"0886",	x"0886",	
												x"08b9",	x"0891",	x"08bc",	x"08a2",	
												x"08bf",	x"08b1",	x"08aa",	x"08b2",	
												x"08d1",	x"08d2",	x"08bb",	x"08b5",	
												x"06d0",	x"0893",	x"0004",	x"000a",	
												x"91d0",	x"7d06",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"1363",	
												x"06cc",	x"06d8",	x"06f8",	x"06de",	
												x"06b9",	x"0704",	x"06e2",	x"06ba",	
												x"06ff",	x"06f7",	x"0711",	x"0704",	
												x"06f0",	x"0701",	x"06e8",	x"06fb",	
												x"06ea",	x"06fa",	x"072d",	x"073c",	
												x"0723",	x"0727",	x"0726",	x"0712",	
												x"0722",	x"0738",	x"072d",	x"0727",	
												x"072c",	x"0739",	x"06ee",	x"073f",	
												x"0709",	x"06fa",	x"0724",	x"071f",	
												x"0719",	x"071b",	x"0736",	x"0730",	
												x"073e",	x"0724",	x"0730",	x"0730",	
												x"0708",	x"0718",	x"06d6",	x"0717",	
												x"0704",	x"0720",	x"071d",	x"071b",	
												x"0738",	x"070d",	x"071b",	x"0721",	
												x"0747",	x"073a",	x"074e",	x"0733",	
												x"071c",	x"0741",	x"06d4",	x"071c",	
												x"102e",	x"1363",	x"06d2",	x"06d5",	
												x"06cc",	x"06dc",	x"06c7",	x"06db",	
												x"06c7",	x"06d3",	x"06fa",	x"06c0",	
												x"06f6",	x"06f6",	x"0710",	x"06f9",	
												x"06d2",	x"0709",	x"0701",	x"0708",	
												x"0707",	x"0703",	x"0711",	x"071d",	
												x"0732",	x"0731",	x"06fa",	x"073e",	
												x"071c",	x"0708",	x"070d",	x"072a",	
												x"06c5",	x"0726",	x"070a",	x"06f9",	
												x"06ff",	x"071d",	x"0712",	x"0710",	
												x"0719",	x"072e",	x"070e",	x"0718",	
												x"06fa",	x"071c",	x"072c",	x"0717",	
												x"06cd",	x"0728",	x"0727",	x"0705",	
												x"0729",	x"0721",	x"0735",	x"071b",	
												x"0723",	x"0722",	x"0739",	x"0737",	
												x"073c",	x"0763",	x"0727",	x"0737",	
												x"06b8",	x"071a",	x"202e",	x"1363",	
												x"06d0",	x"06bf",	x"06cb",	x"06d4",	
												x"06b6",	x"06df",	x"06b6",	x"0697",	
												x"06c0",	x"06cb",	x"06d6",	x"06db",	
												x"06dd",	x"06f5",	x"06bb",	x"06fc",	
												x"06f8",	x"06f2",	x"070a",	x"0710",	
												x"070a",	x"070f",	x"06fe",	x"0711",	
												x"0715",	x"0707",	x"06f8",	x"070b",	
												x"0701",	x"06fc",	x"06c2",	x"070e",	
												x"06cf",	x"06d8",	x"06f6",	x"06da",	
												x"0706",	x"070c",	x"0709",	x"070a",	
												x"0717",	x"06f5",	x"071b",	x"070b",	
												x"070d",	x"06ee",	x"06e2",	x"070d",	
												x"06e8",	x"06fc",	x"0710",	x"06fe",	
												x"071b",	x"0714",	x"071f",	x"071e",	
												x"0720",	x"071d",	x"0728",	x"0728",	
												x"0712",	x"0713",	x"06ad",	x"06e8",	
												x"302e",	x"1363",	x"06be",	x"0685",	
												x"06bf",	x"0693",	x"069e",	x"06ab",	
												x"06dc",	x"06a4",	x"06cb",	x"06c2",	
												x"06e2",	x"06d9",	x"06d6",	x"06e9",	
												x"06c3",	x"06c9",	x"06c1",	x"06c5",	
												x"06e5",	x"06cb",	x"0708",	x"06ef",	
												x"06fb",	x"06f7",	x"06e4",	x"06fc",	
												x"0707",	x"06eb",	x"06e1",	x"070e",	
												x"06c7",	x"06d4",	x"06d3",	x"06c7",	
												x"06f7",	x"06e7",	x"0702",	x"06f8",	
												x"070a",	x"06f7",	x"0714",	x"06fb",	
												x"070b",	x"06ff",	x"06ef",	x"0711",	
												x"06ec",	x"06f2",	x"06e7",	x"06f5",	
												x"0701",	x"06ef",	x"070e",	x"06f6",	
												x"0727",	x"06f6",	x"0723",	x"06f4",	
												x"0724",	x"0708",	x"0726",	x"0709",	
												x"06d7",	x"06f9",	x"0004",	x"000a",	
												x"1dae",	x"51c9",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"1364",	
												x"06d2",	x"06c9",	x"06e6",	x"06a5",	
												x"06e6",	x"06d2",	x"06da",	x"06d9",	
												x"06ea",	x"06cd",	x"06e8",	x"06e0",	
												x"0701",	x"0701",	x"06e0",	x"071d",	
												x"06f9",	x"06d8",	x"0701",	x"0710",	
												x"0711",	x"0716",	x"0728",	x"0707",	
												x"0721",	x"071c",	x"0728",	x"0733",	
												x"0728",	x"071d",	x"06cb",	x"072c",	
												x"071c",	x"070e",	x"070e",	x"0714",	
												x"0738",	x"070f",	x"0746",	x"0748",	
												x"0734",	x"0741",	x"0737",	x"072c",	
												x"0737",	x"0748",	x"0728",	x"072a",	
												x"0740",	x"0743",	x"0746",	x"074d",	
												x"0756",	x"074c",	x"0753",	x"074c",	
												x"0763",	x"0752",	x"0784",	x"0761",	
												x"077a",	x"0752",	x"0703",	x"0747",	
												x"502e",	x"1364",	x"0710",	x"06db",	
												x"0733",	x"0708",	x"06f7",	x"0706",	
												x"0712",	x"070d",	x"0715",	x"070e",	
												x"0750",	x"06fd",	x"0749",	x"0738",	
												x"0727",	x"0736",	x"074a",	x"0720",	
												x"075a",	x"074b",	x"074a",	x"074b",	
												x"0763",	x"075d",	x"075e",	x"0755",	
												x"076a",	x"0750",	x"073d",	x"0751",	
												x"072e",	x"071b",	x"073c",	x"0735",	
												x"0766",	x"072f",	x"0769",	x"0738",	
												x"0783",	x"0773",	x"0780",	x"0750",	
												x"0778",	x"0761",	x"0785",	x"075f",	
												x"073d",	x"0745",	x"0770",	x"074e",	
												x"07a2",	x"0765",	x"078e",	x"0773",	
												x"0796",	x"0771",	x"07a0",	x"076b",	
												x"079b",	x"0783",	x"078f",	x"0782",	
												x"0716",	x"0763",	x"602e",	x"1364",	
												x"071e",	x"06dc",	x"072e",	x"071b",	
												x"0719",	x"06fd",	x"0731",	x"0716",	
												x"0757",	x"072b",	x"0754",	x"0733",	
												x"0755",	x"0740",	x"072d",	x"072b",	
												x"076b",	x"0716",	x"07ad",	x"0777",	
												x"077a",	x"0784",	x"078a",	x"0785",	
												x"079f",	x"0781",	x"0784",	x"0793",	
												x"077f",	x"076d",	x"0770",	x"075f",	
												x"078f",	x"0752",	x"0794",	x"079b",	
												x"07ab",	x"078c",	x"07d4",	x"07a5",	
												x"07c2",	x"07ae",	x"07ad",	x"079b",	
												x"0799",	x"079a",	x"0793",	x"0796",	
												x"07c3",	x"0797",	x"07c2",	x"07cd",	
												x"07d8",	x"079b",	x"07ef",	x"07c2",	
												x"07e5",	x"07bc",	x"07f2",	x"07c0",	
												x"07cd",	x"07ba",	x"0736",	x"07a1",	
												x"702e",	x"1364",	x"0757",	x"0725",	
												x"0768",	x"076c",	x"0758",	x"0753",	
												x"0795",	x"0751",	x"0781",	x"0752",	
												x"07b8",	x"077e",	x"07a7",	x"07c1",	
												x"0755",	x"07ae",	x"07ca",	x"0760",	
												x"07e7",	x"07d1",	x"07f7",	x"07d4",	
												x"0822",	x"080e",	x"07f1",	x"07ed",	
												x"07eb",	x"07f7",	x"07ea",	x"07ca",	
												x"07be",	x"07de",	x"07d8",	x"07b1",	
												x"07ed",	x"07c3",	x"0822",	x"07ce",	
												x"0823",	x"0808",	x"0836",	x"0804",	
												x"083c",	x"081d",	x"080a",	x"080f",	
												x"0815",	x"081f",	x"0826",	x"083c",	
												x"082c",	x"0805",	x"083e",	x"0819",	
												x"087a",	x"0836",	x"0868",	x"0831",	
												x"0875",	x"083f",	x"0842",	x"0852",	
												x"0731",	x"083d",	x"0004",	x"000a",	
												x"5cae",	x"86e1",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"2365",	
												x"075a",	x"073c",	x"0766",	x"0755",	
												x"0786",	x"079c",	x"0788",	x"0778",	
												x"07a5",	x"078c",	x"0798",	x"07bc",	
												x"078c",	x"07a6",	x"0782",	x"079a",	
												x"07a4",	x"0783",	x"07b0",	x"07b8",	
												x"07a2",	x"07c7",	x"07a1",	x"07cf",	
												x"07a7",	x"079f",	x"07a2",	x"07a8",	
												x"0753",	x"07a9",	x"076b",	x"078d",	
												x"078a",	x"0783",	x"078c",	x"079b",	
												x"079b",	x"0797",	x"079c",	x"07b6",	
												x"078a",	x"07d0",	x"07cc",	x"0796",	
												x"07b6",	x"07dc",	x"077f",	x"0798",	
												x"079e",	x"07ab",	x"078f",	x"0786",	
												x"079d",	x"07d5",	x"07cb",	x"079b",	
												x"07d0",	x"07a1",	x"07bb",	x"07c9",	
												x"07b7",	x"0795",	x"0746",	x"07bd",	
												x"102e",	x"2365",	x"0752",	x"074b",	
												x"073e",	x"0752",	x"0760",	x"0758",	
												x"0751",	x"078d",	x"0778",	x"0778",	
												x"077a",	x"0763",	x"077b",	x"0788",	
												x"074e",	x"0788",	x"079b",	x"0784",	
												x"07c1",	x"07ae",	x"07a0",	x"07b8",	
												x"0769",	x"079f",	x"0767",	x"0798",	
												x"0787",	x"0797",	x"0756",	x"07a7",	
												x"0754",	x"07a1",	x"0776",	x"0775",	
												x"0777",	x"0794",	x"0791",	x"0789",	
												x"0777",	x"0792",	x"0778",	x"0787",	
												x"0795",	x"079f",	x"07a6",	x"078e",	
												x"0749",	x"07bb",	x"078b",	x"07a0",	
												x"079b",	x"0794",	x"07ac",	x"07ab",	
												x"0779",	x"07a1",	x"07ac",	x"07bb",	
												x"07bc",	x"07ad",	x"07a3",	x"07b5",	
												x"0741",	x"079b",	x"202e",	x"2365",	
												x"0748",	x"0743",	x"0720",	x"0728",	
												x"0713",	x"073a",	x"071b",	x"0741",	
												x"0754",	x"0761",	x"0765",	x"0783",	
												x"075b",	x"0786",	x"0759",	x"0779",	
												x"075c",	x"0763",	x"0761",	x"077a",	
												x"0772",	x"076a",	x"0770",	x"0775",	
												x"0777",	x"0781",	x"0775",	x"078f",	
												x"0770",	x"078a",	x"072e",	x"076a",	
												x"0779",	x"072e",	x"0777",	x"0775",	
												x"0776",	x"0769",	x"075d",	x"0780",	
												x"0764",	x"0768",	x"0770",	x"077e",	
												x"074e",	x"076e",	x"073a",	x"0756",	
												x"0784",	x"076a",	x"0774",	x"0769",	
												x"0771",	x"0769",	x"076b",	x"0770",	
												x"0780",	x"0772",	x"078c",	x"078b",	
												x"079e",	x"077d",	x"06ea",	x"0789",	
												x"302e",	x"2365",	x"0708",	x"06fb",	
												x"073a",	x"0709",	x"073b",	x"070a",	
												x"0735",	x"073b",	x"072d",	x"0757",	
												x"0735",	x"073b",	x"0731",	x"072b",	
												x"071e",	x"072c",	x"075e",	x"073a",	
												x"076c",	x"0745",	x"075b",	x"076c",	
												x"0773",	x"0767",	x"0763",	x"0759",	
												x"074c",	x"077b",	x"076a",	x"075d",	
												x"0716",	x"0751",	x"0736",	x"0728",	
												x"0756",	x"0753",	x"0772",	x"0758",	
												x"0774",	x"074b",	x"076b",	x"0753",	
												x"0771",	x"0764",	x"0765",	x"0753",	
												x"0750",	x"0750",	x"077a",	x"074e",	
												x"0775",	x"0751",	x"0775",	x"0769",	
												x"0798",	x"0768",	x"079a",	x"0771",	
												x"0783",	x"076c",	x"079c",	x"0764",	
												x"0718",	x"076c",	x"0004",	x"000a",	
												x"586e",	x"cee1",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"2366",	
												x"0729",	x"070a",	x"0751",	x"0724",	
												x"0745",	x"0736",	x"073e",	x"073c",	
												x"073e",	x"075b",	x"0752",	x"0759",	
												x"0737",	x"0735",	x"0744",	x"0754",	
												x"0759",	x"0759",	x"0774",	x"0776",	
												x"077c",	x"0781",	x"077f",	x"07a0",	
												x"076f",	x"0780",	x"0775",	x"0779",	
												x"0770",	x"0789",	x"076e",	x"077c",	
												x"076b",	x"077b",	x"0773",	x"0782",	
												x"0768",	x"0796",	x"07b9",	x"07b5",	
												x"07b2",	x"07a4",	x"079a",	x"07b1",	
												x"079d",	x"07b2",	x"0796",	x"07b2",	
												x"0797",	x"07b6",	x"0796",	x"07a6",	
												x"079c",	x"07a2",	x"07b5",	x"07a3",	
												x"07c1",	x"07ca",	x"07bb",	x"07d3",	
												x"07b7",	x"07c4",	x"0735",	x"07c6",	
												x"502e",	x"2366",	x"075f",	x"0726",	
												x"0768",	x"0770",	x"0768",	x"0770",	
												x"0798",	x"0772",	x"078f",	x"077e",	
												x"07b2",	x"079c",	x"07a2",	x"07af",	
												x"07b1",	x"07b9",	x"07cd",	x"07b3",	
												x"07d1",	x"07c5",	x"07c8",	x"07ce",	
												x"07b6",	x"07d2",	x"07cc",	x"07bf",	
												x"07c1",	x"07b4",	x"07ba",	x"07b3",	
												x"0796",	x"07bd",	x"07c3",	x"0792",	
												x"07c6",	x"07ba",	x"07d1",	x"07a2",	
												x"0813",	x"07b7",	x"0805",	x"07ba",	
												x"07d5",	x"07d1",	x"07e3",	x"07d0",	
												x"07d3",	x"07da",	x"07d5",	x"07df",	
												x"07f2",	x"07a9",	x"07fa",	x"07dc",	
												x"0808",	x"07e7",	x"0814",	x"07d6",	
												x"080c",	x"07ee",	x"0808",	x"07e3",	
												x"074c",	x"07da",	x"602e",	x"2366",	
												x"076e",	x"073a",	x"07b9",	x"075e",	
												x"077b",	x"0781",	x"0791",	x"0781",	
												x"07a4",	x"0790",	x"07ad",	x"079d",	
												x"078d",	x"07bc",	x"07c7",	x"07a4",	
												x"07fe",	x"07d9",	x"07f3",	x"07f6",	
												x"07f3",	x"07e3",	x"0804",	x"07f4",	
												x"0807",	x"07e4",	x"0806",	x"07f8",	
												x"07e8",	x"07e9",	x"07d3",	x"07c8",	
												x"07d6",	x"07b0",	x"07fb",	x"07e9",	
												x"080b",	x"07e2",	x"0815",	x"07fc",	
												x"0818",	x"07ee",	x"0809",	x"080c",	
												x"0815",	x"0809",	x"0802",	x"0804",	
												x"082f",	x"0810",	x"0823",	x"0817",	
												x"0840",	x"0810",	x"0864",	x"0824",	
												x"085b",	x"0822",	x"0853",	x"0822",	
												x"0834",	x"0822",	x"07c4",	x"0815",	
												x"702e",	x"2366",	x"07ba",	x"0771",	
												x"07da",	x"07ad",	x"07cc",	x"07b5",	
												x"07f2",	x"07c6",	x"0816",	x"07d3",	
												x"083c",	x"0816",	x"07ce",	x"082f",	
												x"07fb",	x"07ee",	x"0877",	x"081f",	
												x"085c",	x"0849",	x"083a",	x"0852",	
												x"0850",	x"0822",	x"0852",	x"0839",	
												x"0868",	x"0848",	x"0831",	x"0832",	
												x"083f",	x"0831",	x"085c",	x"0834",	
												x"0879",	x"0858",	x"0868",	x"085f",	
												x"0884",	x"085c",	x"0871",	x"0861",	
												x"0886",	x"0892",	x"087a",	x"087f",	
												x"0869",	x"085b",	x"0888",	x"0894",	
												x"08a6",	x"0892",	x"08a7",	x"087c",	
												x"08f9",	x"0886",	x"08da",	x"087a",	
												x"08db",	x"08a5",	x"08bd",	x"08c9",	
												x"06e7",	x"0898",	x"0004",	x"000a",	
												x"8f1b",	x"fc80",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002e",	x"3367",	
												x"069e",	x"06e3",	x"06ab",	x"06a8",	
												x"06b2",	x"06c9",	x"06fe",	x"06ab",	
												x"06d1",	x"06f4",	x"06f3",	x"06ff",	
												x"06d9",	x"070a",	x"06eb",	x"06f6",	
												x"06e0",	x"06e1",	x"06f8",	x"071f",	
												x"0702",	x"071d",	x"0729",	x"074f",	
												x"06f6",	x"0726",	x"06f4",	x"0710",	
												x"06c7",	x"070a",	x"06e4",	x"06d6",	
												x"06ff",	x"06ec",	x"06fc",	x"070a",	
												x"06fc",	x"0712",	x"06ff",	x"0703",	
												x"0707",	x"0709",	x"06ff",	x"070f",	
												x"071a",	x"06f5",	x"06f9",	x"0721",	
												x"06d5",	x"071b",	x"0724",	x"06f9",	
												x"06f6",	x"0719",	x"06eb",	x"070f",	
												x"06f6",	x"06fc",	x"0720",	x"071f",	
												x"071e",	x"06fb",	x"06c8",	x"06ff",	
												x"102e",	x"3367",	x"06b7",	x"06bb",	
												x"06ab",	x"06d4",	x"0695",	x"06c4",	
												x"06cb",	x"06c6",	x"06e1",	x"06d0",	
												x"06e0",	x"06db",	x"06e4",	x"06da",	
												x"06d6",	x"06ec",	x"070a",	x"06f0",	
												x"0731",	x"06fe",	x"0707",	x"0726",	
												x"06f3",	x"0701",	x"06d9",	x"0708",	
												x"06d2",	x"06e4",	x"06ba",	x"06eb",	
												x"06d1",	x"06ba",	x"06e1",	x"06e1",	
												x"06dc",	x"0704",	x"06f5",	x"0708",	
												x"06f4",	x"070b",	x"06f8",	x"070e",	
												x"0718",	x"0720",	x"06ea",	x"071e",	
												x"06d3",	x"06f9",	x"0703",	x"06e3",	
												x"06fa",	x"0708",	x"070a",	x"06f7",	
												x"06eb",	x"0710",	x"0706",	x"06f3",	
												x"072a",	x"0707",	x"071f",	x"0719",	
												x"069d",	x"0718",	x"202e",	x"3367",	
												x"0687",	x"0694",	x"06a6",	x"06a0",	
												x"06bf",	x"06b8",	x"06b4",	x"06c3",	
												x"06c2",	x"06bb",	x"06bb",	x"06da",	
												x"06a9",	x"06d2",	x"06c5",	x"06db",	
												x"06f4",	x"06e4",	x"06ef",	x"070e",	
												x"06f1",	x"0701",	x"06e2",	x"06f2",	
												x"06dd",	x"06f0",	x"06d8",	x"06e4",	
												x"06c7",	x"06bf",	x"06ab",	x"06d1",	
												x"06e8",	x"06b4",	x"06cf",	x"06dd",	
												x"06d8",	x"06df",	x"06d0",	x"06e6",	
												x"06c4",	x"06de",	x"06d5",	x"06c7",	
												x"06e5",	x"06d1",	x"06dc",	x"06ed",	
												x"06e2",	x"06fd",	x"06fb",	x"06f2",	
												x"06d6",	x"06f9",	x"06f8",	x"06df",	
												x"06dd",	x"0705",	x"06fa",	x"06dd",	
												x"0708",	x"06e1",	x"06a3",	x"06e9",	
												x"302e",	x"3367",	x"06ac",	x"068f",	
												x"0696",	x"06aa",	x"066a",	x"06a5",	
												x"06b2",	x"068b",	x"06a3",	x"0690",	
												x"06da",	x"06d2",	x"06a0",	x"06c2",	
												x"068c",	x"069d",	x"06d4",	x"06a2",	
												x"06c2",	x"06cd",	x"06d4",	x"06c0",	
												x"06cb",	x"06cd",	x"06c4",	x"06d0",	
												x"06c5",	x"06b7",	x"06db",	x"06b2",	
												x"06a1",	x"06c3",	x"06dd",	x"06a7",	
												x"06d6",	x"06dc",	x"06e8",	x"06e2",	
												x"06f0",	x"0713",	x"06de",	x"06d8",	
												x"06fc",	x"06f1",	x"06da",	x"06dc",	
												x"06d5",	x"06cd",	x"06f8",	x"06ce",	
												x"06e5",	x"06e9",	x"06ff",	x"06b0",	
												x"06f8",	x"06eb",	x"0706",	x"06df",	
												x"070b",	x"06e8",	x"070b",	x"06e6",	
												x"06a5",	x"06e3",	x"0004",	x"000a",	
												x"0ec3",	x"c467",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402e",	x"3368",	
												x"06ae",	x"0688",	x"06b1",	x"069d",	
												x"06cf",	x"06a9",	x"06cd",	x"06c6",	
												x"06ac",	x"06bc",	x"06c4",	x"06ac",	
												x"06d4",	x"06b4",	x"06cf",	x"06d8",	
												x"06dd",	x"06d7",	x"06fc",	x"0703",	
												x"06f6",	x"06fa",	x"06f8",	x"0700",	
												x"06f7",	x"06f1",	x"06e0",	x"070a",	
												x"06e4",	x"06fd",	x"06d4",	x"06f1",	
												x"06f1",	x"06f8",	x"06f9",	x"06f1",	
												x"0707",	x"0719",	x"0703",	x"0716",	
												x"0715",	x"0715",	x"070d",	x"0718",	
												x"0731",	x"0714",	x"070e",	x"0727",	
												x"0712",	x"070d",	x"070c",	x"0726",	
												x"072c",	x"0710",	x"073a",	x"072f",	
												x"073a",	x"072f",	x"073a",	x"072f",	
												x"074b",	x"073c",	x"06cc",	x"072d",	
												x"502e",	x"3368",	x"06cf",	x"06d8",	
												x"06e0",	x"06be",	x"06e7",	x"06ad",	
												x"06ea",	x"06d2",	x"06f3",	x"06e1",	
												x"0709",	x"06cd",	x"0719",	x"06fc",	
												x"06fb",	x"0718",	x"072f",	x"06f2",	
												x"0727",	x"072b",	x"0729",	x"0743",	
												x"071b",	x"0743",	x"071d",	x"0726",	
												x"071c",	x"0722",	x"0709",	x"0718",	
												x"06fb",	x"0711",	x"0723",	x"070d",	
												x"0731",	x"071f",	x"072c",	x"071d",	
												x"0738",	x"0720",	x"0749",	x"0729",	
												x"0749",	x"0716",	x"073f",	x"0727",	
												x"074a",	x"0713",	x"075f",	x"072b",	
												x"0752",	x"072d",	x"0766",	x"072f",	
												x"0765",	x"0737",	x"075d",	x"0740",	
												x"0771",	x"0745",	x"0769",	x"0740",	
												x"06c4",	x"074a",	x"602e",	x"3368",	
												x"06e0",	x"06bd",	x"06f1",	x"06be",	
												x"06fa",	x"06e0",	x"0703",	x"06ed",	
												x"06ec",	x"06f0",	x"073c",	x"06e7",	
												x"0715",	x"0726",	x"0721",	x"0707",	
												x"0741",	x"0702",	x"075f",	x"0742",	
												x"074a",	x"072e",	x"0759",	x"072f",	
												x"074c",	x"0757",	x"0754",	x"0737",	
												x"0746",	x"0745",	x"071f",	x"074f",	
												x"076a",	x"0720",	x"0748",	x"0756",	
												x"0761",	x"074f",	x"0780",	x"074e",	
												x"0774",	x"0760",	x"0777",	x"0784",	
												x"077d",	x"0766",	x"076c",	x"0767",	
												x"0770",	x"077e",	x"079e",	x"0776",	
												x"078c",	x"0778",	x"07a6",	x"0768",	
												x"07a8",	x"0779",	x"07aa",	x"077f",	
												x"07b9",	x"0789",	x"0717",	x"076a",	
												x"702e",	x"3368",	x"074d",	x"071d",	
												x"0724",	x"072d",	x"072a",	x"0738",	
												x"074e",	x"0721",	x"071c",	x"072b",	
												x"0760",	x"0731",	x"0763",	x"0754",	
												x"077a",	x"0750",	x"07aa",	x"077b",	
												x"07cf",	x"079e",	x"0790",	x"07a5",	
												x"07ce",	x"077e",	x"07c2",	x"07b1",	
												x"07f3",	x"07ac",	x"0791",	x"0788",	
												x"079a",	x"07a3",	x"07c4",	x"07b3",	
												x"07d6",	x"079c",	x"07cb",	x"07ac",	
												x"07f4",	x"07c4",	x"07d2",	x"07dc",	
												x"07ee",	x"07dc",	x"07f1",	x"07dc",	
												x"07a5",	x"07cc",	x"07de",	x"07ab",	
												x"07de",	x"07e3",	x"0830",	x"07e8",	
												x"0836",	x"07f0",	x"0830",	x"07da",	
												x"082c",	x"081e",	x"081b",	x"0822",	
												x"079c",	x"0813",	x"0004",	x"000a",	
												x"4427",	x"eed3",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"0369",	
												x"0790",	x"078a",	x"0792",	x"07a7",	
												x"0792",	x"077e",	x"07bc",	x"0784",	
												x"0762",	x"0793",	x"0762",	x"0762",	
												x"076f",	x"076e",	x"0766",	x"078b",	
												x"078f",	x"0791",	x"07a2",	x"07a1",	
												x"07c0",	x"07ba",	x"07af",	x"07c6",	
												x"07b0",	x"07c9",	x"07d2",	x"07da",	
												x"07bf",	x"07c2",	x"078b",	x"07ca",	
												x"078f",	x"078d",	x"079c",	x"07a2",	
												x"07a5",	x"07b8",	x"07a5",	x"079e",	
												x"079a",	x"07b0",	x"079b",	x"07a2",	
												x"078a",	x"07a9",	x"077f",	x"07af",	
												x"07c8",	x"07ae",	x"07b2",	x"07bf",	
												x"07ba",	x"079a",	x"07b1",	x"07bf",	
												x"07c4",	x"07b3",	x"07bf",	x"07bb",	
												x"07c3",	x"07b1",	x"0771",	x"07a1",	
												x"102f",	x"0369",	x"077d",	x"0794",	
												x"0775",	x"0772",	x"0769",	x"079f",	
												x"074c",	x"075a",	x"074e",	x"0741",	
												x"0724",	x"0749",	x"0735",	x"0749",	
												x"075e",	x"075c",	x"078e",	x"077c",	
												x"079c",	x"0797",	x"07bc",	x"07ab",	
												x"0798",	x"07ac",	x"0790",	x"07a5",	
												x"0787",	x"07b7",	x"0783",	x"078a",	
												x"0775",	x"078b",	x"078f",	x"078b",	
												x"07b4",	x"07aa",	x"079f",	x"07bf",	
												x"07bc",	x"078e",	x"0781",	x"07a4",	
												x"079f",	x"078d",	x"07ad",	x"0781",	
												x"076e",	x"079c",	x"079d",	x"079d",	
												x"07a4",	x"07c9",	x"07b6",	x"07ae",	
												x"079f",	x"07cb",	x"07de",	x"07a7",	
												x"07d0",	x"07ca",	x"07b9",	x"07bd",	
												x"0784",	x"079c",	x"202f",	x"0369",	
												x"0764",	x"075f",	x"075d",	x"0777",	
												x"0757",	x"077f",	x"073a",	x"0755",	
												x"075d",	x"0752",	x"0749",	x"0750",	
												x"0758",	x"0742",	x"0756",	x"0776",	
												x"077c",	x"075e",	x"0775",	x"079c",	
												x"077a",	x"077b",	x"0777",	x"07a6",	
												x"0789",	x"078e",	x"075e",	x"0779",	
												x"076c",	x"0761",	x"0737",	x"0764",	
												x"0759",	x"076c",	x"0781",	x"0765",	
												x"0792",	x"0780",	x"078b",	x"079c",	
												x"076c",	x"077f",	x"0792",	x"0778",	
												x"07a2",	x"078c",	x"0779",	x"0795",	
												x"078a",	x"0785",	x"0785",	x"0783",	
												x"078b",	x"077d",	x"07ac",	x"07a7",	
												x"079d",	x"0798",	x"079a",	x"079c",	
												x"0797",	x"0776",	x"0758",	x"07ab",	
												x"302f",	x"0369",	x"074e",	x"0756",	
												x"074d",	x"0745",	x"0763",	x"0755",	
												x"076b",	x"0756",	x"0754",	x"0743",	
												x"0761",	x"0732",	x"0750",	x"074e",	
												x"0745",	x"074d",	x"077c",	x"0732",	
												x"078b",	x"0765",	x"0794",	x"074f",	
												x"078e",	x"0776",	x"0797",	x"0782",	
												x"0787",	x"0796",	x"0786",	x"0781",	
												x"0746",	x"0772",	x"079e",	x"0751",	
												x"0792",	x"078a",	x"07a2",	x"0777",	
												x"078e",	x"0785",	x"07a2",	x"0767",	
												x"07b9",	x"0790",	x"07b1",	x"0798",	
												x"078b",	x"0783",	x"07b3",	x"0777",	
												x"079c",	x"0784",	x"07c4",	x"0764",	
												x"07ca",	x"07a6",	x"07b5",	x"07a3",	
												x"07cf",	x"0799",	x"07dc",	x"07a4",	
												x"0794",	x"07a7",	x"0004",	x"000a",	
												x"650b",	x"566f",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"036a",	
												x"078f",	x"076d",	x"076a",	x"0787",	
												x"0774",	x"0765",	x"0780",	x"0746",	
												x"0765",	x"0743",	x"079e",	x"0779",	
												x"0783",	x"07a2",	x"078e",	x"075d",	
												x"0786",	x"0757",	x"07b3",	x"076f",	
												x"07c5",	x"0792",	x"07c8",	x"07af",	
												x"07c7",	x"07a8",	x"07c2",	x"07ba",	
												x"07bb",	x"07ae",	x"07b6",	x"07a2",	
												x"07c8",	x"07c9",	x"07e9",	x"07c7",	
												x"07ce",	x"07cf",	x"07fc",	x"07ce",	
												x"07fb",	x"07d6",	x"07f7",	x"07d2",	
												x"0801",	x"07c4",	x"0804",	x"07d5",	
												x"0804",	x"07c5",	x"0825",	x"07e5",	
												x"082b",	x"07f0",	x"0821",	x"0802",	
												x"0814",	x"07ef",	x"0844",	x"07fa",	
												x"084d",	x"07f8",	x"07f6",	x"080d",	
												x"502f",	x"036a",	x"079f",	x"0790",	
												x"07a7",	x"07a3",	x"07c8",	x"079b",	
												x"07c6",	x"07bf",	x"07c8",	x"0788",	
												x"07c6",	x"07c5",	x"07ea",	x"0781",	
												x"07ff",	x"07d5",	x"07f3",	x"07cc",	
												x"07e5",	x"07f4",	x"0809",	x"07fa",	
												x"07ff",	x"0808",	x"0802",	x"07d2",	
												x"080c",	x"07f1",	x"080f",	x"07f1",	
												x"07eb",	x"07f1",	x"0809",	x"07bc",	
												x"07f0",	x"07db",	x"0804",	x"07b6",	
												x"0810",	x"07d4",	x"0817",	x"07d6",	
												x"083f",	x"07f6",	x"082f",	x"07f3",	
												x"0806",	x"07f7",	x"087d",	x"07e7",	
												x"0853",	x"0815",	x"0860",	x"080e",	
												x"0887",	x"081d",	x"0868",	x"0811",	
												x"0861",	x"082a",	x"0858",	x"0811",	
												x"07fe",	x"0822",	x"602f",	x"036a",	
												x"07df",	x"07cc",	x"0815",	x"07b2",	
												x"07d9",	x"07bf",	x"07fc",	x"07ae",	
												x"07e4",	x"07b4",	x"07c7",	x"07bf",	
												x"081d",	x"07b0",	x"0829",	x"07ce",	
												x"0812",	x"07dd",	x"083a",	x"07ed",	
												x"0821",	x"07ef",	x"0818",	x"07d2",	
												x"0820",	x"07fc",	x"0833",	x"07f6",	
												x"083a",	x"07f2",	x"0844",	x"07f6",	
												x"0838",	x"07f3",	x"0855",	x"080c",	
												x"0832",	x"0819",	x"085e",	x"082b",	
												x"0867",	x"0814",	x"085d",	x"0817",	
												x"086d",	x"0813",	x"0864",	x"081e",	
												x"0871",	x"082d",	x"088b",	x"0822",	
												x"089d",	x"083e",	x"08b6",	x"0864",	
												x"08bb",	x"084d",	x"08b3",	x"0853",	
												x"08af",	x"0870",	x"07f0",	x"0881",	
												x"702f",	x"036a",	x"0828",	x"07b5",	
												x"0800",	x"07de",	x"0803",	x"07af",	
												x"081e",	x"07b9",	x"07e9",	x"077c",	
												x"081d",	x"0790",	x"0815",	x"07b8",	
												x"0800",	x"07fb",	x"0857",	x"07fb",	
												x"084a",	x"0820",	x"0886",	x"0830",	
												x"088b",	x"0867",	x"08ad",	x"0864",	
												x"08aa",	x"0872",	x"0892",	x"0857",	
												x"0876",	x"0864",	x"08ba",	x"0839",	
												x"08cc",	x"0866",	x"08c3",	x"085d",	
												x"08d1",	x"0878",	x"08ed",	x"0885",	
												x"08e2",	x"08ce",	x"08bb",	x"086f",	
												x"08ca",	x"088f",	x"08c8",	x"08a7",	
												x"0909",	x"088f",	x"0905",	x"08a3",	
												x"08fd",	x"0901",	x"08f6",	x"08bc",	
												x"0927",	x"08c3",	x"090d",	x"08db",	
												x"06f9",	x"08e8",	x"0004",	x"000a",	
												x"b473",	x"8de6",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"136b",	
												x"0711",	x"070d",	x"0717",	x"0721",	
												x"06f0",	x"0712",	x"0709",	x"06fa",	
												x"06ec",	x"06e3",	x"06f1",	x"06f8",	
												x"06bd",	x"06e0",	x"06d3",	x"06d9",	
												x"06db",	x"06d5",	x"071c",	x"06f8",	
												x"0724",	x"0720",	x"06f8",	x"0736",	
												x"0734",	x"0722",	x"0755",	x"0743",	
												x"06ff",	x"075b",	x"06ed",	x"071b",	
												x"0718",	x"071b",	x"072f",	x"072e",	
												x"0719",	x"0727",	x"0723",	x"073a",	
												x"072e",	x"0733",	x"0729",	x"074b",	
												x"071b",	x"072e",	x"06f3",	x"0730",	
												x"0721",	x"0703",	x"073d",	x"0741",	
												x"0740",	x"0739",	x"0710",	x"072c",	
												x"0740",	x"0720",	x"0745",	x"0727",	
												x"071d",	x"0738",	x"0705",	x"0715",	
												x"102f",	x"136b",	x"06c9",	x"06c8",	
												x"06ca",	x"06e0",	x"06c5",	x"06ee",	
												x"06d0",	x"06dd",	x"06d1",	x"06ca",	
												x"06c5",	x"06c2",	x"06d6",	x"06d1",	
												x"06a6",	x"06af",	x"0708",	x"06b9",	
												x"070e",	x"071a",	x"06ec",	x"0705",	
												x"0728",	x"072c",	x"0716",	x"073b",	
												x"0713",	x"0729",	x"0709",	x"072b",	
												x"06ed",	x"0718",	x"0706",	x"06fd",	
												x"071e",	x"0707",	x"071c",	x"0732",	
												x"071c",	x"071a",	x"0718",	x"071e",	
												x"072b",	x"071d",	x"0724",	x"072b",	
												x"06e8",	x"0711",	x"0724",	x"0708",	
												x"0734",	x"0713",	x"0744",	x"0727",	
												x"072b",	x"0750",	x"073c",	x"073c",	
												x"0759",	x"072e",	x"0738",	x"0747",	
												x"06e3",	x"0734",	x"202f",	x"136b",	
												x"06fb",	x"06e7",	x"06e2",	x"06fb",	
												x"06f3",	x"06f1",	x"06de",	x"0706",	
												x"06d5",	x"06a1",	x"06df",	x"06f6",	
												x"06af",	x"070a",	x"06ba",	x"06ee",	
												x"06c0",	x"06ef",	x"06f0",	x"06fa",	
												x"0719",	x"0719",	x"0714",	x"0713",	
												x"06f5",	x"071d",	x"06f1",	x"06f4",	
												x"0723",	x"0703",	x"06e0",	x"070b",	
												x"06ee",	x"06f1",	x"06dd",	x"0703",	
												x"0709",	x"06fd",	x"071d",	x"070f",	
												x"0713",	x"06f9",	x"0709",	x"070b",	
												x"0717",	x"0701",	x"06d5",	x"0706",	
												x"06f9",	x"071f",	x"0723",	x"0714",	
												x"0712",	x"071b",	x"0714",	x"0715",	
												x"0720",	x"06f3",	x"071d",	x"072d",	
												x"0720",	x"0706",	x"06d2",	x"06f7",	
												x"302f",	x"136b",	x"06d5",	x"06bf",	
												x"06e3",	x"06be",	x"06c0",	x"06cc",	
												x"06bb",	x"06c0",	x"06e9",	x"06a9",	
												x"06b8",	x"06ae",	x"06aa",	x"06b8",	
												x"06a1",	x"06b0",	x"06de",	x"06ac",	
												x"06ef",	x"06d3",	x"071d",	x"06e4",	
												x"0719",	x"0700",	x"070d",	x"06d1",	
												x"070d",	x"0713",	x"06f5",	x"06ed",	
												x"06ee",	x"06df",	x"0709",	x"06e6",	
												x"070a",	x"06fe",	x"070f",	x"070d",	
												x"0733",	x"070d",	x"072d",	x"071e",	
												x"0718",	x"0702",	x"0726",	x"0700",	
												x"06f2",	x"071c",	x"070e",	x"06f9",	
												x"0747",	x"06f4",	x"0746",	x"070d",	
												x"0747",	x"0714",	x"0743",	x"071a",	
												x"073a",	x"071e",	x"0739",	x"0717",	
												x"06e4",	x"071a",	x"0004",	x"000a",	
												x"21d8",	x"5445",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"136c",	
												x"06c9",	x"06ad",	x"06f4",	x"06c9",	
												x"06fc",	x"06d0",	x"0702",	x"06f8",	
												x"06f9",	x"06d6",	x"06d4",	x"06db",	
												x"06e1",	x"06d1",	x"06ef",	x"06f1",	
												x"0749",	x"06e2",	x"0739",	x"0715",	
												x"072f",	x"0725",	x"0731",	x"0727",	
												x"0739",	x"0720",	x"0743",	x"073f",	
												x"074a",	x"071e",	x"072d",	x"0748",	
												x"073b",	x"0718",	x"0752",	x"0742",	
												x"0756",	x"074e",	x"0767",	x"074d",	
												x"073c",	x"0751",	x"0759",	x"0742",	
												x"0743",	x"0748",	x"074c",	x"0735",	
												x"0796",	x"074e",	x"076e",	x"076e",	
												x"0761",	x"0754",	x"0773",	x"075b",	
												x"0784",	x"0765",	x"0792",	x"0775",	
												x"0782",	x"0768",	x"073b",	x"0730",	
												x"502f",	x"136c",	x"0731",	x"06ff",	
												x"0715",	x"0715",	x"071a",	x"06da",	
												x"0712",	x"0700",	x"0730",	x"06f0",	
												x"0752",	x"06fd",	x"0744",	x"06e2",	
												x"0707",	x"0718",	x"0782",	x"0713",	
												x"0761",	x"074f",	x"0779",	x"073a",	
												x"0775",	x"0756",	x"0767",	x"0768",	
												x"0775",	x"075c",	x"076a",	x"0756",	
												x"0749",	x"0746",	x"0787",	x"073e",	
												x"0795",	x"0765",	x"0792",	x"0771",	
												x"07ac",	x"077a",	x"07a6",	x"0768",	
												x"0795",	x"077b",	x"078d",	x"075b",	
												x"0796",	x"075d",	x"07b3",	x"078e",	
												x"07d0",	x"0793",	x"07b9",	x"0785",	
												x"07ad",	x"0793",	x"07d8",	x"078b",	
												x"07cb",	x"0794",	x"079b",	x"078e",	
												x"073a",	x"0764",	x"602f",	x"136c",	
												x"074a",	x"06f8",	x"074d",	x"0724",	
												x"0739",	x"0732",	x"074e",	x"071b",	
												x"0769",	x"071d",	x"0757",	x"06f8",	
												x"075b",	x"074e",	x"074d",	x"0727",	
												x"076e",	x"0712",	x"0777",	x"077d",	
												x"0780",	x"0772",	x"07ad",	x"0780",	
												x"07b4",	x"077f",	x"07b2",	x"0788",	
												x"07a6",	x"0786",	x"07a2",	x"0793",	
												x"07b8",	x"0785",	x"07ca",	x"079e",	
												x"07fd",	x"07a9",	x"07cb",	x"07b1",	
												x"07d3",	x"07a7",	x"07d8",	x"0799",	
												x"07cd",	x"079d",	x"07c0",	x"07af",	
												x"07e1",	x"07a3",	x"07f0",	x"07b7",	
												x"07f3",	x"07a5",	x"07fe",	x"07b0",	
												x"07ec",	x"07c4",	x"07f4",	x"07d3",	
												x"07d7",	x"07bd",	x"075c",	x"07b2",	
												x"702f",	x"136c",	x"0779",	x"0712",	
												x"07bc",	x"076f",	x"0775",	x"076b",	
												x"07a4",	x"0750",	x"0797",	x"0726",	
												x"0783",	x"074c",	x"0781",	x"0741",	
												x"07bd",	x"0755",	x"07b7",	x"0779",	
												x"07e0",	x"079a",	x"07f8",	x"07b2",	
												x"082a",	x"07ec",	x"081d",	x"07ee",	
												x"0830",	x"0801",	x"082c",	x"07ec",	
												x"07ff",	x"07bf",	x"0827",	x"07bd",	
												x"086b",	x"080d",	x"083f",	x"081a",	
												x"0832",	x"0811",	x"0846",	x"0816",	
												x"0856",	x"080e",	x"081c",	x"0821",	
												x"080d",	x"084d",	x"084f",	x"0823",	
												x"0881",	x"084b",	x"0879",	x"080a",	
												x"0870",	x"0841",	x"088d",	x"0830",	
												x"08a9",	x"0851",	x"0856",	x"0845",	
												x"0763",	x"081c",	x"0004",	x"000a",	
												x"6b7a",	x"89d8",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"236d",	
												x"0774",	x"075a",	x"078d",	x"075d",	
												x"0761",	x"078f",	x"078b",	x"0770",	
												x"075e",	x"0764",	x"0787",	x"075a",	
												x"0776",	x"076c",	x"0782",	x"0784",	
												x"07b9",	x"078a",	x"07c6",	x"07b7",	
												x"07cb",	x"07c8",	x"07b0",	x"07c1",	
												x"07a4",	x"07af",	x"079b",	x"07a4",	
												x"07a3",	x"0794",	x"0769",	x"07a0",	
												x"07ac",	x"0783",	x"07a7",	x"07ca",	
												x"07be",	x"07b5",	x"079c",	x"07bd",	
												x"07a9",	x"07a5",	x"078b",	x"0798",	
												x"07bb",	x"07ad",	x"07bb",	x"079d",	
												x"0798",	x"07cc",	x"07b7",	x"07b6",	
												x"07d7",	x"07bc",	x"07cd",	x"07be",	
												x"07a3",	x"0797",	x"07dd",	x"07b3",	
												x"0796",	x"079a",	x"0765",	x"0789",	
												x"102f",	x"236d",	x"0757",	x"0768",	
												x"0752",	x"0755",	x"0740",	x"076b",	
												x"0720",	x"073f",	x"076f",	x"0749",	
												x"075c",	x"0768",	x"0755",	x"076f",	
												x"075b",	x"0769",	x"079d",	x"0744",	
												x"07a4",	x"079e",	x"078f",	x"0799",	
												x"0781",	x"079e",	x"0784",	x"078e",	
												x"0788",	x"0790",	x"078a",	x"07af",	
												x"0747",	x"07bf",	x"076a",	x"075c",	
												x"07a5",	x"07aa",	x"078b",	x"07b1",	
												x"0799",	x"07a9",	x"0794",	x"07b6",	
												x"07a6",	x"07b5",	x"0792",	x"07ac",	
												x"0757",	x"079b",	x"078d",	x"07b9",	
												x"07a5",	x"07ae",	x"07b2",	x"07bc",	
												x"07a1",	x"07a3",	x"07ab",	x"07ab",	
												x"07c9",	x"079e",	x"07a0",	x"079d",	
												x"0708",	x"07bc",	x"202f",	x"236d",	
												x"0727",	x"071f",	x"0746",	x"0730",	
												x"0753",	x"076c",	x"0745",	x"0763",	
												x"0732",	x"073b",	x"0762",	x"0741",	
												x"0768",	x"0779",	x"0726",	x"0766",	
												x"076b",	x"073a",	x"0780",	x"078e",	
												x"0770",	x"077a",	x"0767",	x"0787",	
												x"0784",	x"078d",	x"078b",	x"0784",	
												x"07a5",	x"0783",	x"076f",	x"0773",	
												x"0782",	x"076e",	x"0787",	x"0786",	
												x"0785",	x"0752",	x"0768",	x"0786",	
												x"078d",	x"0778",	x"0789",	x"0790",	
												x"0797",	x"0798",	x"0787",	x"0786",	
												x"0787",	x"0784",	x"077d",	x"0782",	
												x"0790",	x"0787",	x"0773",	x"079c",	
												x"078c",	x"0786",	x"07d3",	x"0782",	
												x"0793",	x"0790",	x"0737",	x"0771",	
												x"302f",	x"236d",	x"0723",	x"071d",	
												x"0732",	x"0725",	x"072c",	x"0728",	
												x"072f",	x"073d",	x"0721",	x"0713",	
												x"074a",	x"072e",	x"0755",	x"0728",	
												x"0718",	x"0734",	x"0747",	x"0747",	
												x"0753",	x"0758",	x"0769",	x"075d",	
												x"0769",	x"076c",	x"073f",	x"0751",	
												x"074c",	x"0747",	x"0751",	x"0766",	
												x"073e",	x"075a",	x"076f",	x"0745",	
												x"0766",	x"0763",	x"0778",	x"0766",	
												x"076e",	x"075f",	x"0779",	x"075e",	
												x"079b",	x"0767",	x"0777",	x"0761",	
												x"0771",	x"0760",	x"07ce",	x"0764",	
												x"0795",	x"0767",	x"078d",	x"0770",	
												x"0794",	x"0769",	x"07a4",	x"075f",	
												x"0799",	x"077c",	x"0796",	x"077e",	
												x"0734",	x"0769",	x"0004",	x"000a",	
												x"5dcb",	x"cfe0",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"236e",	
												x"0757",	x"0722",	x"0731",	x"0741",	
												x"0747",	x"071a",	x"075c",	x"073b",	
												x"075c",	x"073e",	x"0763",	x"0756",	
												x"0763",	x"0747",	x"076d",	x"0757",	
												x"0785",	x"074f",	x"0785",	x"078d",	
												x"078f",	x"078b",	x"079a",	x"0790",	
												x"0796",	x"078a",	x"078d",	x"0794",	
												x"079b",	x"0797",	x"079f",	x"078c",	
												x"07c5",	x"079d",	x"07b3",	x"07c3",	
												x"07cf",	x"07b0",	x"07ca",	x"079b",	
												x"07c3",	x"07a2",	x"07bd",	x"07d0",	
												x"07b5",	x"07cf",	x"07b7",	x"07c5",	
												x"07d1",	x"07c9",	x"07cf",	x"07bf",	
												x"07d4",	x"07c9",	x"07c0",	x"07e0",	
												x"07e9",	x"07d0",	x"07df",	x"07d8",	
												x"07c9",	x"07cb",	x"0769",	x"07c0",	
												x"502f",	x"236e",	x"076a",	x"073b",	
												x"0777",	x"0762",	x"079b",	x"0737",	
												x"07a8",	x"077f",	x"07a8",	x"0776",	
												x"077d",	x"0783",	x"07d6",	x"0774",	
												x"07ac",	x"07c3",	x"07b9",	x"0794",	
												x"07e1",	x"07b4",	x"07d0",	x"07c8",	
												x"07e2",	x"07c0",	x"0805",	x"07b6",	
												x"07dd",	x"07c9",	x"07da",	x"07c7",	
												x"07e3",	x"07b8",	x"07ff",	x"07b9",	
												x"0801",	x"07d8",	x"07f6",	x"07b8",	
												x"081b",	x"07d9",	x"0821",	x"07e9",	
												x"080f",	x"07fb",	x"0842",	x"07f1",	
												x"0803",	x"0807",	x"081f",	x"07fe",	
												x"0818",	x"07dc",	x"0826",	x"07dd",	
												x"083d",	x"07de",	x"0849",	x"07d7",	
												x"083d",	x"07fb",	x"0821",	x"07ff",	
												x"077f",	x"07e8",	x"602f",	x"236e",	
												x"0784",	x"0772",	x"07c8",	x"0769",	
												x"0799",	x"0780",	x"07ab",	x"078a",	
												x"07cb",	x"075c",	x"07da",	x"0766",	
												x"07e5",	x"07b6",	x"0802",	x"07c4",	
												x"082b",	x"07bd",	x"0829",	x"07cc",	
												x"0829",	x"07e8",	x"0852",	x"0803",	
												x"081b",	x"07eb",	x"0825",	x"07f6",	
												x"0829",	x"07f1",	x"0809",	x"07d9",	
												x"0847",	x"07ea",	x"0828",	x"080e",	
												x"0833",	x"07e9",	x"0853",	x"07fe",	
												x"085a",	x"0812",	x"0846",	x"0813",	
												x"0866",	x"0818",	x"0849",	x"080c",	
												x"083d",	x"082a",	x"0837",	x"081e",	
												x"0867",	x"0818",	x"0873",	x"082f",	
												x"0873",	x"0831",	x"087c",	x"0829",	
												x"0862",	x"083d",	x"07e6",	x"0813",	
												x"702f",	x"236e",	x"07e0",	x"0780",	
												x"07da",	x"079d",	x"07e8",	x"0789",	
												x"07fe",	x"07a1",	x"07f8",	x"07c6",	
												x"082c",	x"07ea",	x"0842",	x"07d3",	
												x"07f3",	x"07f7",	x"084c",	x"07d0",	
												x"086d",	x"0817",	x"088b",	x"082d",	
												x"0895",	x"084f",	x"08b6",	x"082c",	
												x"08a1",	x"0863",	x"0878",	x"085f",	
												x"087d",	x"083c",	x"087c",	x"083d",	
												x"088d",	x"084f",	x"0881",	x"085a",	
												x"08c3",	x"0885",	x"08ba",	x"0899",	
												x"08cf",	x"088b",	x"08c3",	x"0897",	
												x"0894",	x"08ab",	x"08a9",	x"088e",	
												x"08bb",	x"08b6",	x"08b1",	x"08b3",	
												x"08ec",	x"08b7",	x"08f0",	x"0890",	
												x"08f6",	x"08bf",	x"08d6",	x"08ae",	
												x"0703",	x"08d3",	x"0004",	x"000a",	
												x"a23a",	x"00ba",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"002f",	x"336f",	
												x"06da",	x"06ec",	x"06dd",	x"06f8",	
												x"06cf",	x"06ce",	x"06c9",	x"06dc",	
												x"06f3",	x"06cb",	x"06ff",	x"06fc",	
												x"06af",	x"06d7",	x"06f2",	x"06ca",	
												x"070d",	x"06d5",	x"06f8",	x"0727",	
												x"06fc",	x"071f",	x"0720",	x"0727",	
												x"0707",	x"0739",	x"071a",	x"073c",	
												x"06fb",	x"0730",	x"06d7",	x"06f4",	
												x"071c",	x"06fc",	x"06e6",	x"06f2",	
												x"06fd",	x"0705",	x"0701",	x"0709",	
												x"0707",	x"070b",	x"071c",	x"071e",	
												x"070f",	x"0727",	x"06d9",	x"0721",	
												x"0708",	x"070d",	x"0723",	x"071c",	
												x"06f9",	x"0723",	x"06e6",	x"06f9",	
												x"06e7",	x"0706",	x"0704",	x"0717",	
												x"06f7",	x"0700",	x"06bc",	x"06f9",	
												x"102f",	x"336f",	x"06cc",	x"06c9",	
												x"06bd",	x"06bf",	x"06bb",	x"06c3",	
												x"06bb",	x"06ce",	x"06b8",	x"06bd",	
												x"06c2",	x"06b4",	x"06c8",	x"06c6",	
												x"069a",	x"06c5",	x"0702",	x"06c9",	
												x"0728",	x"06fe",	x"06fd",	x"0707",	
												x"06ee",	x"0704",	x"06fb",	x"0702",	
												x"0700",	x"06e0",	x"06ff",	x"06f8",	
												x"06e1",	x"06f2",	x"06fa",	x"06c9",	
												x"06ef",	x"070a",	x"06ee",	x"070e",	
												x"06eb",	x"06e4",	x"06d3",	x"06f8",	
												x"070b",	x"06f7",	x"0714",	x"0711",	
												x"06ef",	x"0705",	x"0725",	x"06fb",	
												x"0700",	x"0725",	x"06fe",	x"0713",	
												x"06e7",	x"0718",	x"0708",	x"06fd",	
												x"071a",	x"0719",	x"0720",	x"070a",	
												x"06c2",	x"0725",	x"202f",	x"336f",	
												x"06b6",	x"06b3",	x"06ae",	x"06b6",	
												x"06c6",	x"068a",	x"0690",	x"06b0",	
												x"0681",	x"0699",	x"0690",	x"06a9",	
												x"0681",	x"06a3",	x"06b1",	x"06b7",	
												x"06e1",	x"06cc",	x"06e9",	x"06f3",	
												x"06e7",	x"06f7",	x"06f1",	x"06e6",	
												x"06d6",	x"06ec",	x"06de",	x"06fe",	
												x"06e9",	x"06bf",	x"06bf",	x"06df",	
												x"0702",	x"06d1",	x"06e3",	x"06f9",	
												x"06eb",	x"06e0",	x"06e7",	x"06f3",	
												x"06dd",	x"06e3",	x"06e8",	x"06e4",	
												x"06e3",	x"06f7",	x"06cc",	x"06ea",	
												x"06e6",	x"06f0",	x"06e2",	x"06ee",	
												x"06fb",	x"06ef",	x"06f1",	x"06f3",	
												x"06e3",	x"06e3",	x"0707",	x"06f4",	
												x"0704",	x"06f1",	x"06ca",	x"06ea",	
												x"302f",	x"336f",	x"06b1",	x"069b",	
												x"06b0",	x"069d",	x"0680",	x"0688",	
												x"06a6",	x"0685",	x"0697",	x"0683",	
												x"0695",	x"068e",	x"06b2",	x"06a4",	
												x"06ab",	x"06a9",	x"06d4",	x"06bb",	
												x"06e0",	x"06c4",	x"06da",	x"06c3",	
												x"06df",	x"06d1",	x"06e8",	x"06d3",	
												x"06e6",	x"06c8",	x"06e1",	x"06c2",	
												x"06d0",	x"06d3",	x"06ce",	x"06b2",	
												x"06d7",	x"06e4",	x"06f1",	x"06e2",	
												x"070e",	x"0708",	x"06e3",	x"06fb",	
												x"0709",	x"06f2",	x"070e",	x"06d8",	
												x"06f3",	x"06ce",	x"0708",	x"06d4",	
												x"070f",	x"0710",	x"0714",	x"06f1",	
												x"0704",	x"06d8",	x"0710",	x"06d8",	
												x"0703",	x"06de",	x"06f3",	x"06de",	
												x"06b1",	x"06d7",	x"0004",	x"000a",	
												x"11c2",	x"c47c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"402f",	x"3370",	
												x"06b8",	x"0684",	x"06b3",	x"06a1",	
												x"06ce",	x"0680",	x"06d1",	x"06af",	
												x"06cb",	x"06ac",	x"06d3",	x"06a7",	
												x"06e8",	x"06ae",	x"06ed",	x"06b9",	
												x"06f9",	x"06ef",	x"070e",	x"06ee",	
												x"06ef",	x"06ec",	x"06e6",	x"06ee",	
												x"0704",	x"06e1",	x"0709",	x"06ed",	
												x"0723",	x"0715",	x"06e5",	x"0711",	
												x"0725",	x"070d",	x"072a",	x"0708",	
												x"0727",	x"0736",	x"0721",	x"0728",	
												x"0731",	x"070d",	x"072c",	x"0725",	
												x"0743",	x"0728",	x"0740",	x"0737",	
												x"075f",	x"072d",	x"0742",	x"0738",	
												x"0744",	x"0737",	x"0749",	x"0736",	
												x"0785",	x"073b",	x"0742",	x"0740",	
												x"0749",	x"0738",	x"0702",	x"072a",	
												x"502f",	x"3370",	x"0705",	x"06df",	
												x"0703",	x"06fb",	x"06e2",	x"06ba",	
												x"071d",	x"06e6",	x"0710",	x"0703",	
												x"072d",	x"06df",	x"0720",	x"0706",	
												x"0712",	x"06f4",	x"0731",	x"070f",	
												x"0740",	x"0728",	x"074f",	x"0739",	
												x"074f",	x"0758",	x"0758",	x"073e",	
												x"0754",	x"0738",	x"073f",	x"071c",	
												x"0723",	x"073f",	x"0745",	x"0714",	
												x"0756",	x"0732",	x"0758",	x"073a",	
												x"0772",	x"073f",	x"077c",	x"073c",	
												x"0785",	x"072f",	x"0789",	x"0752",	
												x"075c",	x"0753",	x"07ab",	x"0741",	
												x"075d",	x"075b",	x"0781",	x"0738",	
												x"0787",	x"074a",	x"0793",	x"073e",	
												x"07ab",	x"0764",	x"077a",	x"0763",	
												x"0712",	x"074f",	x"602f",	x"3370",	
												x"0729",	x"06f7",	x"0721",	x"06f1",	
												x"06e5",	x"06d5",	x"073a",	x"06db",	
												x"071b",	x"06ec",	x"0732",	x"0700",	
												x"0736",	x"071e",	x"0739",	x"0727",	
												x"0761",	x"071b",	x"077a",	x"0746",	
												x"077c",	x"075a",	x"078e",	x"074e",	
												x"077c",	x"0772",	x"0780",	x"0761",	
												x"0778",	x"0772",	x"0770",	x"074b",	
												x"0791",	x"0738",	x"079a",	x"0789",	
												x"0784",	x"0779",	x"0798",	x"0778",	
												x"0789",	x"0786",	x"07a6",	x"077e",	
												x"07a4",	x"076f",	x"07a4",	x"07a2",	
												x"07bb",	x"077b",	x"07bb",	x"07a0",	
												x"07c5",	x"0778",	x"07b9",	x"077c",	
												x"07c5",	x"077b",	x"07ac",	x"078d",	
												x"07b4",	x"0795",	x"072b",	x"077a",	
												x"702f",	x"3370",	x"0746",	x"0701",	
												x"0743",	x"0707",	x"0742",	x"0702",	
												x"0751",	x"0700",	x"075c",	x"0718",	
												x"075f",	x"0727",	x"07a1",	x"0742",	
												x"0775",	x"075e",	x"07aa",	x"0769",	
												x"07d4",	x"079b",	x"07ca",	x"0781",	
												x"07df",	x"078f",	x"07e5",	x"0788",	
												x"07ce",	x"07ab",	x"07db",	x"07a1",	
												x"07ab",	x"07bd",	x"07f7",	x"0777",	
												x"0814",	x"07c9",	x"07c4",	x"07b3",	
												x"07d0",	x"07bb",	x"07d7",	x"07c4",	
												x"0823",	x"07ca",	x"0833",	x"07de",	
												x"07ef",	x"07dd",	x"083a",	x"07e7",	
												x"083c",	x"07f5",	x"0835",	x"07d9",	
												x"0820",	x"07d2",	x"0854",	x"07ea",	
												x"0854",	x"07fa",	x"0823",	x"0817",	
												x"0787",	x"07ff",	x"0004",	x"000a",	
												x"548a",	x"f3a1",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"0371",	
												x"0799",	x"07d1",	x"0785",	x"07ba",	
												x"0786",	x"0793",	x"07a8",	x"076e",	
												x"07a9",	x"07b2",	x"07e2",	x"07ee",	
												x"07d7",	x"07f8",	x"07b5",	x"07e6",	
												x"07be",	x"07d6",	x"07bd",	x"07a8",	
												x"07bf",	x"0812",	x"07bf",	x"07d9",	
												x"07b4",	x"07d9",	x"07ca",	x"07f9",	
												x"07cd",	x"07dd",	x"077c",	x"07e7",	
												x"078d",	x"07b2",	x"07a9",	x"07de",	
												x"07ab",	x"07db",	x"07da",	x"07d0",	
												x"07d8",	x"07d9",	x"07d1",	x"0819",	
												x"07bc",	x"07e4",	x"0770",	x"07d6",	
												x"07bb",	x"0791",	x"07ff",	x"07c3",	
												x"07d3",	x"07c5",	x"0804",	x"07fe",	
												x"0802",	x"07e1",	x"07ea",	x"07f5",	
												x"07ee",	x"07d8",	x"07a2",	x"07f2",	
												x"1030",	x"0371",	x"07a8",	x"080f",	
												x"07a3",	x"07c4",	x"07a9",	x"07be",	
												x"07bb",	x"07bc",	x"07e8",	x"07aa",	
												x"07df",	x"07f8",	x"07f0",	x"07e5",	
												x"07d2",	x"0808",	x"07da",	x"07ff",	
												x"07da",	x"07ca",	x"07d9",	x"07e9",	
												x"07fe",	x"080a",	x"07ea",	x"080d",	
												x"07d9",	x"07e7",	x"07d7",	x"07d5",	
												x"07c8",	x"07e2",	x"07b6",	x"07b1",	
												x"07d7",	x"07fc",	x"07fc",	x"0813",	
												x"07f2",	x"07f9",	x"07fa",	x"0800",	
												x"07e9",	x"0806",	x"0805",	x"07dc",	
												x"0760",	x"07f4",	x"07c6",	x"07b8",	
												x"07eb",	x"07d2",	x"07f8",	x"07f1",	
												x"07f7",	x"07ff",	x"0811",	x"07f5",	
												x"080d",	x"07fc",	x"07ec",	x"0808",	
												x"07a1",	x"07c7",	x"2030",	x"0371",	
												x"0799",	x"07dc",	x"077d",	x"079a",	
												x"078e",	x"07a8",	x"0782",	x"07c7",	
												x"07db",	x"07ec",	x"07dc",	x"07ea",	
												x"07d8",	x"07e6",	x"07a3",	x"07d9",	
												x"07bd",	x"07cd",	x"07ae",	x"07d0",	
												x"07b1",	x"07c5",	x"07ca",	x"07de",	
												x"07bc",	x"07d8",	x"07ce",	x"07dd",	
												x"07c1",	x"07d5",	x"075b",	x"079f",	
												x"07a8",	x"079d",	x"07b6",	x"07e4",	
												x"07be",	x"079a",	x"07c1",	x"07cf",	
												x"07bf",	x"07bb",	x"07c3",	x"07d0",	
												x"07c6",	x"07bc",	x"0771",	x"07c7",	
												x"07d3",	x"07a1",	x"07d9",	x"07d4",	
												x"07ca",	x"07d8",	x"07e1",	x"07e7",	
												x"07e0",	x"07e3",	x"07c4",	x"07e3",	
												x"07e1",	x"079f",	x"0734",	x"07e4",	
												x"3030",	x"0371",	x"0736",	x"0772",	
												x"0735",	x"0729",	x"0757",	x"073c",	
												x"075b",	x"0762",	x"0756",	x"0739",	
												x"0780",	x"078d",	x"0782",	x"0795",	
												x"0771",	x"079b",	x"0793",	x"0776",	
												x"079c",	x"079e",	x"0795",	x"0789",	
												x"0785",	x"0787",	x"0791",	x"078c",	
												x"078f",	x"0787",	x"0777",	x"0768",	
												x"0742",	x"076c",	x"0782",	x"0772",	
												x"078d",	x"07a6",	x"0794",	x"07a7",	
												x"07a8",	x"078d",	x"07bd",	x"07ab",	
												x"07bd",	x"07a3",	x"079a",	x"07ab",	
												x"0732",	x"075e",	x"07ae",	x"077b",	
												x"07af",	x"0794",	x"07da",	x"07a4",	
												x"07d6",	x"07c4",	x"07b6",	x"07a2",	
												x"07d8",	x"0792",	x"07e0",	x"07ae",	
												x"0781",	x"07a3",	x"0004",	x"000a",	
												x"7aae",	x"7397",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"0372",	
												x"076c",	x"0796",	x"074f",	x"075e",	
												x"075c",	x"0736",	x"0790",	x"076b",	
												x"0780",	x"078d",	x"07a3",	x"07a9",	
												x"0798",	x"07aa",	x"0794",	x"0794",	
												x"07b7",	x"0788",	x"07b6",	x"07aa",	
												x"07be",	x"07cb",	x"07b8",	x"07c6",	
												x"07b7",	x"07bc",	x"07b7",	x"07c8",	
												x"07ac",	x"07ca",	x"079d",	x"07bf",	
												x"07ac",	x"079d",	x"07ab",	x"07c4",	
												x"07db",	x"07ae",	x"07f7",	x"07df",	
												x"0800",	x"07f3",	x"07dd",	x"07e0",	
												x"0791",	x"07cf",	x"0799",	x"0796",	
												x"07cb",	x"07a8",	x"080e",	x"07d9",	
												x"080f",	x"07e1",	x"0821",	x"0812",	
												x"0800",	x"07df",	x"0807",	x"07fa",	
												x"082d",	x"07e4",	x"07da",	x"07ec",	
												x"5030",	x"0372",	x"07a0",	x"07bf",	
												x"079b",	x"07a7",	x"07b7",	x"077c",	
												x"07cc",	x"07a6",	x"07c1",	x"07c1",	
												x"07ef",	x"07e2",	x"07cf",	x"07e8",	
												x"07cd",	x"07e1",	x"07e4",	x"07de",	
												x"07ed",	x"07ff",	x"07ff",	x"07e3",	
												x"07fe",	x"07f6",	x"0826",	x"080d",	
												x"07cb",	x"082b",	x"07d8",	x"07c9",	
												x"07db",	x"07cf",	x"07e3",	x"07d9",	
												x"0808",	x"07dd",	x"0818",	x"07de",	
												x"081c",	x"0810",	x"0827",	x"0801",	
												x"0830",	x"080c",	x"081a",	x"07f7",	
												x"0805",	x"07e0",	x"0821",	x"07e9",	
												x"0822",	x"07f5",	x"0842",	x"0802",	
												x"087a",	x"081d",	x"0849",	x"0829",	
												x"0852",	x"0820",	x"084e",	x"0808",	
												x"07d1",	x"0813",	x"6030",	x"0372",	
												x"07b5",	x"07dd",	x"07dc",	x"07b6",	
												x"07ce",	x"07d9",	x"07e4",	x"07c7",	
												x"082c",	x"07d1",	x"07ff",	x"07fa",	
												x"07f7",	x"0803",	x"07f2",	x"07f2",	
												x"0821",	x"07f1",	x"084d",	x"080b",	
												x"0815",	x"080f",	x"0837",	x"0809",	
												x"082b",	x"0812",	x"083b",	x"084f",	
												x"0822",	x"080c",	x"0804",	x"07f7",	
												x"081f",	x"07ea",	x"0826",	x"081b",	
												x"083a",	x"0808",	x"0855",	x"0843",	
												x"0863",	x"082d",	x"086c",	x"084e",	
												x"085c",	x"083c",	x"0847",	x"0812",	
												x"086b",	x"0807",	x"086b",	x"0854",	
												x"0881",	x"084a",	x"088b",	x"085d",	
												x"08c0",	x"0846",	x"088b",	x"085c",	
												x"0891",	x"086b",	x"082f",	x"0867",	
												x"7030",	x"0372",	x"07f4",	x"081e",	
												x"080d",	x"07de",	x"080d",	x"07c8",	
												x"07ff",	x"07ed",	x"0833",	x"082b",	
												x"088c",	x"0818",	x"0870",	x"087d",	
												x"0842",	x"0865",	x"08bf",	x"0854",	
												x"0886",	x"084b",	x"0885",	x"088d",	
												x"08e5",	x"0875",	x"08bb",	x"089c",	
												x"08ae",	x"0894",	x"0878",	x"08a3",	
												x"086f",	x"089d",	x"08bf",	x"087c",	
												x"08ea",	x"08b5",	x"08dd",	x"08b2",	
												x"08f9",	x"08b2",	x"08e3",	x"08b6",	
												x"08c9",	x"08c6",	x"08cd",	x"089f",	
												x"0894",	x"08a8",	x"08fc",	x"08b3",	
												x"0909",	x"08ff",	x"08e8",	x"08f0",	
												x"08fe",	x"0902",	x"08fb",	x"08fc",	
												x"093c",	x"08fc",	x"092c",	x"090b",	
												x"0708",	x"0901",	x"0004",	x"000a",	
												x"b16c",	x"9b18",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"1373",	
												x"06b8",	x"0711",	x"06f8",	x"06cc",	
												x"06dd",	x"06f6",	x"06fa",	x"06e6",	
												x"0713",	x"06ff",	x"0717",	x"0707",	
												x"071a",	x"0722",	x"06e9",	x"0727",	
												x"06ce",	x"06ec",	x"0724",	x"070e",	
												x"0718",	x"0725",	x"071c",	x"070d",	
												x"0727",	x"0747",	x"0734",	x"0738",	
												x"0720",	x"073c",	x"06d9",	x"073b",	
												x"06f0",	x"06f5",	x"0744",	x"0718",	
												x"0721",	x"0713",	x"071f",	x"0738",	
												x"071e",	x"071a",	x"0726",	x"073a",	
												x"071e",	x"0713",	x"06bc",	x"072d",	
												x"0723",	x"06de",	x"0738",	x"0738",	
												x"0739",	x"0730",	x"071c",	x"070c",	
												x"0735",	x"0724",	x"0752",	x"0713",	
												x"0710",	x"0729",	x"06eb",	x"0705",	
												x"1030",	x"1373",	x"06b7",	x"06fa",	
												x"06d2",	x"06c3",	x"06c7",	x"06d3",	
												x"06f7",	x"06e9",	x"0713",	x"06ee",	
												x"0706",	x"070d",	x"0721",	x"071c",	
												x"0716",	x"0714",	x"0723",	x"072c",	
												x"0712",	x"071e",	x"0718",	x"0730",	
												x"0715",	x"0746",	x"0713",	x"0736",	
												x"071f",	x"0724",	x"071d",	x"071f",	
												x"06b8",	x"0722",	x"06fc",	x"06de",	
												x"0708",	x"0713",	x"071b",	x"071d",	
												x"0721",	x"0723",	x"071b",	x"0717",	
												x"06fd",	x"0718",	x"06ff",	x"06ff",	
												x"06f8",	x"0700",	x"0706",	x"06d7",	
												x"0721",	x"070d",	x"0737",	x"0723",	
												x"0714",	x"0721",	x"073d",	x"0735",	
												x"0744",	x"0737",	x"074c",	x"0731",	
												x"06ca",	x"073a",	x"2030",	x"1373",	
												x"06dc",	x"06ca",	x"06d6",	x"06e7",	
												x"06dc",	x"06dd",	x"06cd",	x"06d3",	
												x"06d4",	x"06c8",	x"06f4",	x"06f6",	
												x"06de",	x"0719",	x"06c3",	x"06ff",	
												x"06cc",	x"06ff",	x"06d7",	x"06f6",	
												x"0712",	x"0717",	x"06e3",	x"0729",	
												x"070c",	x"0705",	x"070f",	x"0708",	
												x"070c",	x"070d",	x"06b8",	x"0706",	
												x"06df",	x"06cc",	x"06fb",	x"06f2",	
												x"0714",	x"06f4",	x"0714",	x"0731",	
												x"070c",	x"0708",	x"0702",	x"06f9",	
												x"0715",	x"0700",	x"06d4",	x"0702",	
												x"0704",	x"06d5",	x"0716",	x"0711",	
												x"071f",	x"0707",	x"071c",	x"0707",	
												x"0722",	x"0724",	x"0722",	x"072f",	
												x"070d",	x"0722",	x"06bf",	x"06fc",	
												x"3030",	x"1373",	x"06b1",	x"06b3",	
												x"06c7",	x"0693",	x"06ac",	x"06e0",	
												x"06e1",	x"06b1",	x"06e5",	x"06e0",	
												x"06f2",	x"06ea",	x"06ec",	x"06ec",	
												x"06c2",	x"06e8",	x"06ee",	x"06e6",	
												x"06f5",	x"06e3",	x"06f9",	x"0705",	
												x"06f0",	x"06ee",	x"06ef",	x"06e7",	
												x"06e5",	x"06f7",	x"06dc",	x"06f2",	
												x"06b3",	x"06d8",	x"06eb",	x"06b4",	
												x"06f9",	x"06e1",	x"06fd",	x"06f4",	
												x"0712",	x"0704",	x"0724",	x"070c",	
												x"071b",	x"0721",	x"0718",	x"0716",	
												x"06e3",	x"0712",	x"0709",	x"06f3",	
												x"0720",	x"0701",	x"0718",	x"0709",	
												x"0728",	x"0702",	x"0732",	x"0709",	
												x"0735",	x"071f",	x"0734",	x"070d",	
												x"06a6",	x"06ff",	x"0004",	x"000a",	
												x"200f",	x"54aa",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"1374",	
												x"06ae",	x"06b5",	x"06db",	x"06b6",	
												x"06df",	x"06bd",	x"06ea",	x"06ea",	
												x"06e3",	x"06e9",	x"070b",	x"06df",	
												x"0714",	x"070b",	x"06df",	x"0713",	
												x"0726",	x"06e1",	x"0727",	x"0726",	
												x"0731",	x"0736",	x"072a",	x"072c",	
												x"072f",	x"0721",	x"0739",	x"073a",	
												x"072c",	x"0729",	x"0704",	x"0735",	
												x"0722",	x"06ff",	x"0721",	x"072b",	
												x"0744",	x"0733",	x"074b",	x"0764",	
												x"0743",	x"0746",	x"074b",	x"0755",	
												x"072a",	x"074d",	x"0713",	x"072a",	
												x"074a",	x"0735",	x"0759",	x"0751",	
												x"074f",	x"075f",	x"0761",	x"0758",	
												x"0760",	x"0764",	x"0776",	x"0763",	
												x"0777",	x"075e",	x"071f",	x"0755",	
												x"5030",	x"1374",	x"0725",	x"0726",	
												x"0738",	x"071b",	x"0703",	x"0714",	
												x"0732",	x"0726",	x"0737",	x"0724",	
												x"0750",	x"072c",	x"0764",	x"073d",	
												x"0715",	x"075c",	x"074e",	x"0732",	
												x"078d",	x"074a",	x"0766",	x"0766",	
												x"075b",	x"075b",	x"0756",	x"0754",	
												x"074d",	x"0750",	x"075e",	x"074c",	
												x"0727",	x"075a",	x"0754",	x"0708",	
												x"0767",	x"0749",	x"077d",	x"074b",	
												x"0797",	x"0775",	x"0787",	x"076d",	
												x"0782",	x"076b",	x"077d",	x"075c",	
												x"0761",	x"0730",	x"077e",	x"0758",	
												x"0792",	x"076d",	x"079c",	x"076d",	
												x"079b",	x"078b",	x"07aa",	x"076a",	
												x"07a8",	x"0790",	x"07a0",	x"078f",	
												x"0716",	x"0776",	x"6030",	x"1374",	
												x"0739",	x"070d",	x"0732",	x"0718",	
												x"0713",	x"0721",	x"0761",	x"06fa",	
												x"075b",	x"071f",	x"075e",	x"0744",	
												x"074f",	x"0748",	x"076a",	x"0726",	
												x"0769",	x"0757",	x"0795",	x"0782",	
												x"0784",	x"0785",	x"0791",	x"0795",	
												x"0796",	x"0780",	x"07a8",	x"0793",	
												x"07b0",	x"0780",	x"0771",	x"0787",	
												x"07a1",	x"075e",	x"07aa",	x"079e",	
												x"07b3",	x"0793",	x"07b4",	x"07a5",	
												x"07d1",	x"07a2",	x"07bb",	x"0794",	
												x"07c6",	x"079c",	x"07a3",	x"07c8",	
												x"07cd",	x"07b7",	x"07d3",	x"07c7",	
												x"07ed",	x"07a7",	x"07fd",	x"07c5",	
												x"07fe",	x"07d0",	x"080f",	x"07c9",	
												x"07d4",	x"07e3",	x"0794",	x"07ac",	
												x"7030",	x"1374",	x"076e",	x"078a",	
												x"07d2",	x"0772",	x"077f",	x"0762",	
												x"07c0",	x"0770",	x"07de",	x"07a9",	
												x"07cf",	x"0797",	x"07df",	x"07c9",	
												x"07cf",	x"07df",	x"0812",	x"07ba",	
												x"080c",	x"07d8",	x"0809",	x"07eb",	
												x"0825",	x"0815",	x"081b",	x"0817",	
												x"082c",	x"0827",	x"07f3",	x"0814",	
												x"0804",	x"07eb",	x"0814",	x"07df",	
												x"0834",	x"0823",	x"084d",	x"081a",	
												x"0840",	x"083d",	x"0843",	x"082b",	
												x"0846",	x"0825",	x"0838",	x"082c",	
												x"080f",	x"084e",	x"0858",	x"0831",	
												x"0854",	x"0855",	x"0889",	x"0850",	
												x"0887",	x"085f",	x"0884",	x"0875",	
												x"088e",	x"085e",	x"0870",	x"0867",	
												x"0776",	x"0844",	x"0004",	x"000a",	
												x"66ec",	x"90d9",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"2375",	
												x"0763",	x"079c",	x"0771",	x"076c",	
												x"0764",	x"076e",	x"0795",	x"0788",	
												x"079e",	x"0798",	x"07d4",	x"07b9",	
												x"07ad",	x"07ca",	x"078e",	x"07b6",	
												x"079e",	x"079e",	x"07c4",	x"07c5",	
												x"07d2",	x"07c1",	x"07c2",	x"07d5",	
												x"0791",	x"07d8",	x"079c",	x"0792",	
												x"07ab",	x"0790",	x"074c",	x"0787",	
												x"0793",	x"0762",	x"0785",	x"07af",	
												x"0798",	x"0783",	x"07a9",	x"07be",	
												x"07ad",	x"07a8",	x"07b3",	x"0797",	
												x"07cf",	x"07d0",	x"0749",	x"07ad",	
												x"07a4",	x"0776",	x"07a1",	x"07af",	
												x"07ad",	x"07aa",	x"07ab",	x"0799",	
												x"07a6",	x"0799",	x"07c6",	x"07b8",	
												x"07d2",	x"07bd",	x"0753",	x"07b9",	
												x"1030",	x"2375",	x"074a",	x"0781",	
												x"0750",	x"0753",	x"07a4",	x"0763",	
												x"0775",	x"07ac",	x"0786",	x"078e",	
												x"0778",	x"077e",	x"0781",	x"07a1",	
												x"0784",	x"0781",	x"07b5",	x"0798",	
												x"07c5",	x"07aa",	x"07a7",	x"07a0",	
												x"078d",	x"079d",	x"0775",	x"079c",	
												x"0774",	x"0790",	x"074d",	x"0792",	
												x"0750",	x"0794",	x"076a",	x"0775",	
												x"07ab",	x"0787",	x"078b",	x"07a8",	
												x"0797",	x"07af",	x"078c",	x"079a",	
												x"0798",	x"079b",	x"0787",	x"0790",	
												x"075e",	x"07b6",	x"078b",	x"0793",	
												x"07ae",	x"079f",	x"07b9",	x"07ac",	
												x"077e",	x"07a7",	x"07a5",	x"07b6",	
												x"07bb",	x"07b1",	x"07b4",	x"07ba",	
												x"0756",	x"07b1",	x"2030",	x"2375",	
												x"0727",	x"078a",	x"073d",	x"0715",	
												x"074f",	x"075e",	x"0784",	x"0789",	
												x"0767",	x"0795",	x"0768",	x"0780",	
												x"0768",	x"0781",	x"0756",	x"0783",	
												x"0768",	x"0780",	x"0780",	x"078f",	
												x"079f",	x"0791",	x"0786",	x"078e",	
												x"0761",	x"0792",	x"0797",	x"0783",	
												x"077e",	x"0796",	x"0756",	x"0763",	
												x"075a",	x"073a",	x"0771",	x"0768",	
												x"0779",	x"0780",	x"0758",	x"0786",	
												x"077f",	x"076f",	x"0779",	x"0780",	
												x"077a",	x"0775",	x"0762",	x"075f",	
												x"076f",	x"0762",	x"076a",	x"076f",	
												x"078e",	x"0783",	x"0774",	x"078b",	
												x"0792",	x"0786",	x"0794",	x"0788",	
												x"0786",	x"0772",	x"0700",	x"075c",	
												x"3030",	x"2375",	x"071b",	x"073c",	
												x"072c",	x"070e",	x"0724",	x"0711",	
												x"0739",	x"0727",	x"072e",	x"0748",	
												x"0741",	x"074d",	x"0743",	x"0748",	
												x"0734",	x"072f",	x"074b",	x"0761",	
												x"076c",	x"0753",	x"076f",	x"0778",	
												x"0771",	x"076a",	x"075f",	x"0753",	
												x"0755",	x"0756",	x"075c",	x"076a",	
												x"0713",	x"0743",	x"0751",	x"0759",	
												x"0765",	x"0758",	x"0764",	x"0753",	
												x"0761",	x"0745",	x"0765",	x"076e",	
												x"0784",	x"0776",	x"0780",	x"0765",	
												x"0738",	x"077a",	x"077d",	x"0730",	
												x"0763",	x"0758",	x"0782",	x"0751",	
												x"078a",	x"077c",	x"079e",	x"0772",	
												x"078d",	x"0777",	x"07a1",	x"077a",	
												x"073a",	x"0783",	x"0004",	x"000a",	
												x"5d19",	x"d312",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"2376",	
												x"0738",	x"0751",	x"0758",	x"073c",	
												x"0729",	x"0749",	x"0742",	x"072c",	
												x"0754",	x"0765",	x"075b",	x"0761",	
												x"0767",	x"0753",	x"0755",	x"0769",	
												x"0784",	x"0769",	x"078d",	x"078e",	
												x"0779",	x"0780",	x"077f",	x"0787",	
												x"077c",	x"0789",	x"078a",	x"079a",	
												x"0773",	x"0795",	x"077d",	x"077f",	
												x"0783",	x"078c",	x"078f",	x"0795",	
												x"078e",	x"07a8",	x"078e",	x"07a1",	
												x"078f",	x"07aa",	x"07ab",	x"07c2",	
												x"07a8",	x"07bc",	x"0781",	x"07b6",	
												x"0784",	x"07a3",	x"07a1",	x"0796",	
												x"07ab",	x"07ba",	x"07ee",	x"07c2",	
												x"07cd",	x"07c4",	x"07be",	x"07c7",	
												x"07b4",	x"07c1",	x"0753",	x"07bd",	
												x"5030",	x"2376",	x"0767",	x"0790",	
												x"0778",	x"0760",	x"0785",	x"0763",	
												x"07a7",	x"0779",	x"07b1",	x"07a7",	
												x"07c1",	x"07b5",	x"07a0",	x"07c0",	
												x"07c1",	x"07c1",	x"07ce",	x"07b7",	
												x"07e0",	x"07ab",	x"07de",	x"07d4",	
												x"07c0",	x"07de",	x"07d3",	x"07bf",	
												x"07c4",	x"07e3",	x"07dd",	x"07b6",	
												x"07b3",	x"07a6",	x"07c3",	x"079c",	
												x"07ec",	x"07d3",	x"07ed",	x"07cf",	
												x"07f3",	x"07dc",	x"07f0",	x"07cb",	
												x"07e4",	x"07d0",	x"07e1",	x"07ce",	
												x"07c1",	x"07b6",	x"07f2",	x"07b1",	
												x"07fe",	x"07d4",	x"07fd",	x"07ec",	
												x"084c",	x"07ea",	x"082d",	x"07db",	
												x"0817",	x"07fe",	x"0803",	x"07ed",	
												x"0796",	x"07de",	x"6030",	x"2376",	
												x"079b",	x"0783",	x"07a8",	x"078e",	
												x"0797",	x"079d",	x"07ed",	x"07ae",	
												x"07b9",	x"07af",	x"07b5",	x"07a7",	
												x"07a7",	x"07a6",	x"07b8",	x"07c7",	
												x"0804",	x"07e1",	x"080b",	x"07ea",	
												x"0800",	x"07f1",	x"0813",	x"080b",	
												x"0810",	x"07ce",	x"080e",	x"07ee",	
												x"0810",	x"07fd",	x"0803",	x"07fa",	
												x"0801",	x"07ef",	x"080d",	x"0804",	
												x"0818",	x"07f6",	x"081d",	x"080e",	
												x"0847",	x"081c",	x"0815",	x"081d",	
												x"082b",	x"0800",	x"0811",	x"0809",	
												x"083e",	x"080e",	x"082d",	x"0828",	
												x"0846",	x"0817",	x"0864",	x"083a",	
												x"0860",	x"0827",	x"0862",	x"0840",	
												x"0853",	x"0818",	x"07ee",	x"0818",	
												x"7030",	x"2376",	x"07bc",	x"07d1",	
												x"07dc",	x"07a1",	x"07dc",	x"07d8",	
												x"0848",	x"07ef",	x"080b",	x"07ee",	
												x"0846",	x"0815",	x"0844",	x"083b",	
												x"0844",	x"081e",	x"0869",	x"0837",	
												x"086f",	x"0857",	x"085d",	x"086a",	
												x"0867",	x"085c",	x"0876",	x"085a",	
												x"0888",	x"0872",	x"0851",	x"0881",	
												x"086a",	x"0854",	x"0882",	x"0859",	
												x"08b1",	x"0880",	x"0888",	x"0890",	
												x"08a0",	x"088a",	x"08a5",	x"087e",	
												x"08e4",	x"08b7",	x"08a6",	x"08a5",	
												x"0885",	x"08aa",	x"08c4",	x"08a2",	
												x"08cf",	x"08c0",	x"08cb",	x"08b1",	
												x"08f3",	x"08c5",	x"08f3",	x"08ce",	
												x"08f5",	x"08e5",	x"08d7",	x"08dd",	
												x"06c7",	x"08d7",	x"0004",	x"000a",	
												x"98f8",	x"06aa",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0030",	x"3377",	
												x"06b0",	x"071b",	x"06be",	x"06b0",	
												x"06c8",	x"06bb",	x"06c3",	x"06d9",	
												x"06d4",	x"0702",	x"0710",	x"0706",	
												x"06e1",	x"071e",	x"06dd",	x"0703",	
												x"06da",	x"06da",	x"0741",	x"0717",	
												x"06e4",	x"074d",	x"06e7",	x"0707",	
												x"06f4",	x"06fc",	x"06ea",	x"0723",	
												x"06b7",	x"06e7",	x"069e",	x"06c7",	
												x"06d8",	x"06d8",	x"06da",	x"06db",	
												x"06da",	x"0704",	x"06fa",	x"0700",	
												x"0710",	x"070d",	x"0704",	x"0738",	
												x"06e3",	x"06f3",	x"06e7",	x"0700",	
												x"071f",	x"06f6",	x"06f4",	x"0733",	
												x"06f3",	x"0704",	x"06e3",	x"06fa",	
												x"06ec",	x"070a",	x"0713",	x"070d",	
												x"0729",	x"0725",	x"068c",	x"071a",	
												x"1030",	x"3377",	x"0697",	x"06a3",	
												x"06cc",	x"069d",	x"0692",	x"06d3",	
												x"06dc",	x"06ad",	x"070c",	x"06d3",	
												x"06db",	x"06fa",	x"06da",	x"06ea",	
												x"06c5",	x"06e2",	x"06f6",	x"06e2",	
												x"070e",	x"06f4",	x"0711",	x"0729",	
												x"070e",	x"0711",	x"06f1",	x"070f",	
												x"06f1",	x"06e6",	x"06bb",	x"06e6",	
												x"06cb",	x"06d2",	x"06c8",	x"06e5",	
												x"06d0",	x"06ee",	x"06d6",	x"0703",	
												x"06f5",	x"06f1",	x"06e6",	x"0714",	
												x"06ff",	x"072a",	x"06ff",	x"06fa",	
												x"06cc",	x"06ef",	x"06ec",	x"06ca",	
												x"06e7",	x"06f4",	x"06ee",	x"06eb",	
												x"0705",	x"06f7",	x"0706",	x"070e",	
												x"0717",	x"0710",	x"0739",	x"06ee",	
												x"068b",	x"0734",	x"2030",	x"3377",	
												x"0693",	x"06bf",	x"06a2",	x"0699",	
												x"06ad",	x"06c8",	x"06ab",	x"06b8",	
												x"06c7",	x"06c7",	x"06bf",	x"06d9",	
												x"06ac",	x"06e6",	x"06c3",	x"06fb",	
												x"06d8",	x"06e7",	x"06c7",	x"06ef",	
												x"06d6",	x"06f7",	x"06e5",	x"06f4",	
												x"06d5",	x"06e4",	x"06d4",	x"06ee",	
												x"06d2",	x"06e7",	x"0693",	x"06ef",	
												x"06ed",	x"06c4",	x"06e1",	x"06e3",	
												x"06e9",	x"06e4",	x"06e4",	x"06e7",	
												x"06d9",	x"06d8",	x"06f5",	x"06cc",	
												x"06bb",	x"06da",	x"06ab",	x"06b8",	
												x"06e7",	x"06c2",	x"06f4",	x"06d1",	
												x"06de",	x"06ee",	x"06e1",	x"06e8",	
												x"06f9",	x"06f8",	x"06fd",	x"06f5",	
												x"0703",	x"06ec",	x"069a",	x"0701",	
												x"3030",	x"3377",	x"0682",	x"06ae",	
												x"068b",	x"069f",	x"06a0",	x"0696",	
												x"06b9",	x"0698",	x"069a",	x"069a",	
												x"06bf",	x"06bb",	x"06ab",	x"06c0",	
												x"06a9",	x"06b8",	x"06cf",	x"06b8",	
												x"06dd",	x"06db",	x"06fa",	x"06c5",	
												x"06df",	x"06e7",	x"06ce",	x"06ca",	
												x"06c8",	x"06bc",	x"06c7",	x"06be",	
												x"069e",	x"06da",	x"06cd",	x"06a1",	
												x"06d5",	x"06d0",	x"06de",	x"06cf",	
												x"06ee",	x"06d9",	x"06f4",	x"06d7",	
												x"06e4",	x"06e8",	x"06f6",	x"06d6",	
												x"06bb",	x"06f4",	x"06bc",	x"06ab",	
												x"0711",	x"06c8",	x"06f2",	x"06d2",	
												x"06f4",	x"06cb",	x"0712",	x"06d1",	
												x"0713",	x"06e6",	x"070e",	x"06fd",	
												x"06c1",	x"06df",	x"0004",	x"000a",	
												x"0d04",	x"c44c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4030",	x"3378",	
												x"06ad",	x"06b6",	x"06c3",	x"0682",	
												x"06d1",	x"06ab",	x"06c4",	x"06cd",	
												x"06be",	x"06aa",	x"06b2",	x"06d6",	
												x"06c9",	x"06b7",	x"06cb",	x"06d4",	
												x"06e9",	x"06ce",	x"06f3",	x"06f1",	
												x"06ef",	x"0708",	x"06d9",	x"0704",	
												x"06f8",	x"06e2",	x"06eb",	x"06fd",	
												x"06e9",	x"06ff",	x"06c1",	x"06f9",	
												x"06fa",	x"06d9",	x"06f9",	x"06e4",	
												x"0716",	x"070f",	x"0714",	x"0720",	
												x"0723",	x"0716",	x"0711",	x"071b",	
												x"070b",	x"0719",	x"06fe",	x"06fe",	
												x"0708",	x"06fd",	x"070c",	x"0705",	
												x"0735",	x"0719",	x"072e",	x"072d",	
												x"0759",	x"0727",	x"0746",	x"0747",	
												x"074f",	x"0742",	x"06f8",	x"0731",	
												x"5030",	x"3378",	x"06fa",	x"0701",	
												x"06ed",	x"06da",	x"06e5",	x"06d0",	
												x"06fc",	x"06e7",	x"06f5",	x"06f6",	
												x"06f5",	x"06e9",	x"073c",	x"0703",	
												x"0705",	x"070b",	x"071b",	x"0712",	
												x"0746",	x"071e",	x"0747",	x"0733",	
												x"0731",	x"073d",	x"072c",	x"0722",	
												x"072c",	x"0727",	x"0726",	x"0725",	
												x"06d1",	x"0715",	x"0727",	x"0706",	
												x"0740",	x"0730",	x"073d",	x"072b",	
												x"074d",	x"073f",	x"074f",	x"0731",	
												x"0758",	x"0725",	x"074f",	x"072d",	
												x"0753",	x"073b",	x"076a",	x"0729",	
												x"075f",	x"072f",	x"0764",	x"0730",	
												x"0775",	x"0741",	x"0778",	x"0741",	
												x"076a",	x"074a",	x"077c",	x"0746",	
												x"0732",	x"0761",	x"6030",	x"3378",	
												x"0716",	x"0728",	x"070a",	x"06f4",	
												x"0714",	x"06f9",	x"074b",	x"070b",	
												x"0730",	x"072f",	x"0720",	x"070f",	
												x"0723",	x"0713",	x"0723",	x"071f",	
												x"075f",	x"06ef",	x"0777",	x"0762",	
												x"0767",	x"0757",	x"076d",	x"074a",	
												x"0762",	x"0757",	x"0778",	x"0761",	
												x"0769",	x"075f",	x"073d",	x"0769",	
												x"076a",	x"072a",	x"076d",	x"075b",	
												x"0793",	x"0770",	x"077f",	x"077a",	
												x"0774",	x"0774",	x"079d",	x"0777",	
												x"0796",	x"0789",	x"0774",	x"0773",	
												x"0797",	x"0779",	x"0796",	x"077e",	
												x"0799",	x"0764",	x"07a9",	x"0776",	
												x"07ae",	x"0780",	x"07d9",	x"0785",	
												x"07b1",	x"078d",	x"076f",	x"0771",	
												x"7030",	x"3378",	x"0762",	x"074c",	
												x"0744",	x"0757",	x"0744",	x"0755",	
												x"076e",	x"072d",	x"074d",	x"073d",	
												x"078a",	x"075c",	x"079e",	x"078a",	
												x"07aa",	x"078f",	x"07c1",	x"07a3",	
												x"07d2",	x"07c3",	x"07cf",	x"07cf",	
												x"07e0",	x"07c8",	x"07dd",	x"07b9",	
												x"07d6",	x"07e1",	x"07d2",	x"07a2",	
												x"07c3",	x"07d0",	x"07c3",	x"07ac",	
												x"07e2",	x"07cd",	x"07fe",	x"07d4",	
												x"07e4",	x"07f7",	x"07f3",	x"07f6",	
												x"080b",	x"07f2",	x"0811",	x"07fd",	
												x"07d8",	x"0813",	x"080e",	x"07d8",	
												x"0828",	x"0804",	x"0811",	x"07fd",	
												x"085d",	x"07dd",	x"084a",	x"07f8",	
												x"0843",	x"083b",	x"0834",	x"0822",	
												x"07a1",	x"0815",	x"0004",	x"000a",	
												x"4ce2",	x"f6ed",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"0379",	
												x"0745",	x"0792",	x"078a",	x"0793",	
												x"074d",	x"0744",	x"074f",	x"0748",	
												x"074f",	x"074c",	x"0760",	x"0755",	
												x"0767",	x"0747",	x"0730",	x"0776",	
												x"0792",	x"0787",	x"0796",	x"078e",	
												x"07a4",	x"079f",	x"0796",	x"07a1",	
												x"0795",	x"07bb",	x"07b5",	x"07b2",	
												x"077b",	x"0791",	x"0761",	x"07b4",	
												x"0775",	x"0776",	x"0780",	x"07a0",	
												x"0794",	x"07a6",	x"079b",	x"079c",	
												x"078d",	x"0799",	x"0789",	x"0796",	
												x"078a",	x"07a1",	x"0765",	x"07aa",	
												x"07a1",	x"0780",	x"07a6",	x"07be",	
												x"07b3",	x"079c",	x"0795",	x"07bb",	
												x"07b8",	x"078f",	x"07a2",	x"07a7",	
												x"07a6",	x"077f",	x"0769",	x"079a",	
												x"1031",	x"0379",	x"0765",	x"0795",	
												x"0753",	x"0753",	x"0745",	x"0752",	
												x"0702",	x"072b",	x"071e",	x"0718",	
												x"0712",	x"0729",	x"0755",	x"0720",	
												x"073d",	x"0756",	x"076b",	x"0762",	
												x"0781",	x"0777",	x"0771",	x"0797",	
												x"0775",	x"0792",	x"0774",	x"078b",	
												x"078b",	x"0780",	x"077f",	x"0782",	
												x"0751",	x"077b",	x"0775",	x"0764",	
												x"077c",	x"078a",	x"078c",	x"0781",	
												x"0789",	x"077a",	x"0770",	x"0798",	
												x"0797",	x"0771",	x"078b",	x"079d",	
												x"0753",	x"079f",	x"078b",	x"0756",	
												x"077b",	x"0799",	x"07b6",	x"0797",	
												x"07a5",	x"07c3",	x"07cd",	x"07a4",	
												x"07a6",	x"07af",	x"07a4",	x"07a8",	
												x"0731",	x"0771",	x"2031",	x"0379",	
												x"0764",	x"0734",	x"075c",	x"0761",	
												x"071a",	x"0748",	x"06ef",	x"0746",	
												x"0722",	x"071f",	x"073c",	x"0714",	
												x"074d",	x"0729",	x"073c",	x"0777",	
												x"0770",	x"075e",	x"077a",	x"0781",	
												x"0776",	x"076f",	x"073a",	x"0789",	
												x"0767",	x"0761",	x"0749",	x"0785",	
												x"0742",	x"074f",	x"0724",	x"0750",	
												x"0793",	x"075f",	x"075e",	x"0783",	
												x"076d",	x"075f",	x"075e",	x"076e",	
												x"0751",	x"0749",	x"077a",	x"0772",	
												x"07a0",	x"075e",	x"0767",	x"078c",	
												x"076d",	x"076c",	x"0779",	x"076d",	
												x"0765",	x"0789",	x"0790",	x"0766",	
												x"0799",	x"075a",	x"078a",	x"0784",	
												x"078b",	x"076c",	x"0715",	x"0784",	
												x"3031",	x"0379",	x"0729",	x"0714",	
												x"073d",	x"0728",	x"072c",	x"0721",	
												x"0738",	x"0707",	x"071f",	x"0725",	
												x"0723",	x"06f9",	x"0761",	x"072c",	
												x"0748",	x"0768",	x"074f",	x"073e",	
												x"0760",	x"075b",	x"076c",	x"0745",	
												x"0760",	x"0750",	x"0770",	x"0754",	
												x"0750",	x"0763",	x"0779",	x"073a",	
												x"0740",	x"0737",	x"0788",	x"074f",	
												x"078d",	x"0783",	x"0789",	x"0787",	
												x"078a",	x"077c",	x"0788",	x"0778",	
												x"078d",	x"0773",	x"0798",	x"0787",	
												x"0780",	x"076d",	x"07a8",	x"075b",	
												x"0784",	x"076a",	x"0792",	x"0762",	
												x"079c",	x"0786",	x"079b",	x"0786",	
												x"07a1",	x"0783",	x"07ae",	x"0750",	
												x"0771",	x"0772",	x"0004",	x"000a",	
												x"572f",	x"497c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"037a",	
												x"075d",	x"074d",	x"0774",	x"0752",	
												x"073a",	x"073c",	x"0773",	x"0722",	
												x"0746",	x"072e",	x"0757",	x"0753",	
												x"0759",	x"0754",	x"0779",	x"074b",	
												x"0793",	x"073f",	x"07a4",	x"0765",	
												x"07ba",	x"0784",	x"0798",	x"079b",	
												x"07ac",	x"078b",	x"07b7",	x"07a1",	
												x"07b9",	x"07a6",	x"0795",	x"079c",	
												x"07c1",	x"079e",	x"07ce",	x"079f",	
												x"07c7",	x"07aa",	x"07d6",	x"07b3",	
												x"07d6",	x"07b8",	x"07cb",	x"07b1",	
												x"07d9",	x"07c4",	x"07e2",	x"07aa",	
												x"07e4",	x"07b7",	x"0818",	x"07d1",	
												x"07f9",	x"07e0",	x"07fa",	x"07eb",	
												x"0815",	x"07d0",	x"07fc",	x"07e7",	
												x"07f4",	x"07cd",	x"079b",	x"07c2",	
												x"5031",	x"037a",	x"079d",	x"077d",	
												x"0787",	x"07a4",	x"0783",	x"076a",	
												x"07a8",	x"0779",	x"0791",	x"0767",	
												x"07ae",	x"078e",	x"07b6",	x"079e",	
												x"07ac",	x"07a8",	x"07f0",	x"07c6",	
												x"07df",	x"07d5",	x"07f2",	x"07d5",	
												x"07e5",	x"07df",	x"07f3",	x"07d4",	
												x"07f7",	x"07d2",	x"0806",	x"07cb",	
												x"07c2",	x"07c7",	x"07f3",	x"07a6",	
												x"07f4",	x"07e0",	x"07f8",	x"07bb",	
												x"07ff",	x"07c2",	x"0836",	x"07d8",	
												x"083c",	x"07e4",	x"0821",	x"07dd",	
												x"07f4",	x"07d0",	x"083d",	x"07ee",	
												x"0826",	x"07f4",	x"0835",	x"07f2",	
												x"0837",	x"0807",	x"082e",	x"07e1",	
												x"0839",	x"0801",	x"081b",	x"07ef",	
												x"0796",	x"07e8",	x"6031",	x"037a",	
												x"07c0",	x"0784",	x"07fc",	x"07b1",	
												x"07a9",	x"07a3",	x"07c1",	x"076e",	
												x"07b5",	x"078d",	x"07ed",	x"07ad",	
												x"07ea",	x"0797",	x"07ec",	x"07e3",	
												x"081e",	x"07c5",	x"0826",	x"07e6",	
												x"0812",	x"07fa",	x"081b",	x"07f4",	
												x"084b",	x"0803",	x"082d",	x"07f9",	
												x"0844",	x"0825",	x"080a",	x"07f1",	
												x"0829",	x"07e5",	x"0815",	x"0820",	
												x"083c",	x"0807",	x"0871",	x"080d",	
												x"0880",	x"083d",	x"0846",	x"0832",	
												x"0877",	x"0811",	x"0819",	x"0819",	
												x"0881",	x"0805",	x"0877",	x"0834",	
												x"087e",	x"0825",	x"0877",	x"0845",	
												x"0882",	x"081e",	x"086d",	x"082d",	
												x"086d",	x"084c",	x"082d",	x"0849",	
												x"7031",	x"037a",	x"080a",	x"082a",	
												x"07ff",	x"07db",	x"0815",	x"07ad",	
												x"080e",	x"07d4",	x"0833",	x"07e0",	
												x"085e",	x"07e3",	x"0851",	x"07f5",	
												x"0851",	x"0820",	x"0892",	x"082d",	
												x"088d",	x"0850",	x"0894",	x"0884",	
												x"0897",	x"0893",	x"08bf",	x"087c",	
												x"08c5",	x"087a",	x"08a5",	x"0862",	
												x"0878",	x"0870",	x"08b2",	x"087b",	
												x"08be",	x"0889",	x"08c1",	x"089b",	
												x"08d3",	x"088b",	x"08f4",	x"0895",	
												x"08f3",	x"08af",	x"08de",	x"08a0",	
												x"08bd",	x"08a3",	x"08f1",	x"08a3",	
												x"092e",	x"08cb",	x"091f",	x"08f6",	
												x"08ff",	x"08e9",	x"0900",	x"08d1",	
												x"0915",	x"08f0",	x"08fd",	x"08be",	
												x"06db",	x"08e9",	x"0004",	x"000a",	
												x"abf8",	x"89f0",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"137b",	
												x"0717",	x"0700",	x"0715",	x"06f2",	
												x"06ed",	x"06f3",	x"06e6",	x"06d7",	
												x"06e8",	x"06dc",	x"06db",	x"06e1",	
												x"06c4",	x"06de",	x"06d6",	x"06cd",	
												x"06fa",	x"06d5",	x"0706",	x"070e",	
												x"0708",	x"0711",	x"06f5",	x"0702",	
												x"070a",	x"0728",	x"0714",	x"072e",	
												x"0709",	x"0729",	x"06d0",	x"0718",	
												x"06e2",	x"071f",	x"072e",	x"070c",	
												x"0713",	x"0709",	x"0717",	x"072c",	
												x"0726",	x"070d",	x"0716",	x"071b",	
												x"0702",	x"06ff",	x"06df",	x"0730",	
												x"06ff",	x"06d9",	x"072f",	x"0714",	
												x"0725",	x"070d",	x"071f",	x"0720",	
												x"0722",	x"06e1",	x"0731",	x"0716",	
												x"06f6",	x"071d",	x"0709",	x"0711",	
												x"1031",	x"137b",	x"06f8",	x"06fd",	
												x"06da",	x"06fa",	x"06c1",	x"06ee",	
												x"06b4",	x"06d2",	x"06c0",	x"0697",	
												x"06e2",	x"06c1",	x"06d1",	x"06cb",	
												x"06b9",	x"06bc",	x"0701",	x"06d0",	
												x"0710",	x"06e7",	x"06f2",	x"06fd",	
												x"06ed",	x"0704",	x"06ff",	x"0705",	
												x"071a",	x"071c",	x"06ec",	x"0706",	
												x"06db",	x"070a",	x"06e9",	x"06fc",	
												x"0720",	x"06e0",	x"0703",	x"0722",	
												x"0703",	x"0709",	x"06ef",	x"0711",	
												x"06f3",	x"0707",	x"06f0",	x"06fd",	
												x"06fc",	x"0700",	x"070e",	x"06ea",	
												x"0715",	x"070f",	x"071c",	x"0709",	
												x"0711",	x"071f",	x"0728",	x"0720",	
												x"072a",	x"0718",	x"073c",	x"0724",	
												x"06bf",	x"0722",	x"2031",	x"137b",	
												x"06d3",	x"06ed",	x"06e6",	x"06e1",	
												x"06c7",	x"06c9",	x"06be",	x"06cf",	
												x"06ad",	x"06cc",	x"06b8",	x"06a4",	
												x"06cc",	x"06c6",	x"06a5",	x"06ec",	
												x"06b9",	x"06e6",	x"06f8",	x"0703",	
												x"0713",	x"0706",	x"0706",	x"070f",	
												x"06f3",	x"06f6",	x"06f3",	x"0709",	
												x"06f2",	x"0704",	x"06b5",	x"06f9",	
												x"06ef",	x"06d4",	x"06e9",	x"06f9",	
												x"06fb",	x"06fc",	x"06f8",	x"0705",	
												x"06fd",	x"06e7",	x"071a",	x"06eb",	
												x"0702",	x"06f8",	x"06eb",	x"0713",	
												x"06f8",	x"06d8",	x"071f",	x"0715",	
												x"0711",	x"0713",	x"0712",	x"0706",	
												x"071f",	x"070e",	x"0728",	x"072a",	
												x"0723",	x"0720",	x"06cf",	x"06e9",	
												x"3031",	x"137b",	x"06c4",	x"06c5",	
												x"06b8",	x"0694",	x"06ca",	x"06a6",	
												x"06cd",	x"06d2",	x"06a2",	x"06af",	
												x"06ad",	x"06ac",	x"0699",	x"06a7",	
												x"0690",	x"069e",	x"06da",	x"0691",	
												x"0702",	x"06d6",	x"0712",	x"06d1",	
												x"070e",	x"06f3",	x"06ec",	x"06e6",	
												x"06fa",	x"06d5",	x"06ec",	x"06e8",	
												x"06e0",	x"06df",	x"06fb",	x"06dc",	
												x"06ff",	x"0701",	x"070a",	x"0703",	
												x"0716",	x"06ff",	x"0712",	x"071b",	
												x"070e",	x"06f2",	x"070e",	x"070f",	
												x"06f4",	x"0704",	x"0707",	x"06e4",	
												x"0729",	x"06e8",	x"0731",	x"0709",	
												x"0750",	x"0701",	x"0734",	x"0709",	
												x"072b",	x"070b",	x"071b",	x"0703",	
												x"06e3",	x"06e8",	x"0004",	x"000a",	
												x"1af8",	x"4c22",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"137c",	
												x"06ec",	x"06d6",	x"06fb",	x"06df",	
												x"06ff",	x"06e2",	x"06ce",	x"06ef",	
												x"06e5",	x"06c1",	x"06e4",	x"06c6",	
												x"06f2",	x"06d0",	x"06f3",	x"06d0",	
												x"0718",	x"06ed",	x"0715",	x"070e",	
												x"073c",	x"0718",	x"071a",	x"0728",	
												x"072b",	x"0723",	x"0740",	x"0737",	
												x"0734",	x"072a",	x"071e",	x"072d",	
												x"0729",	x"071f",	x"0752",	x"072f",	
												x"0757",	x"0740",	x"0756",	x"074e",	
												x"073b",	x"073e",	x"076e",	x"073e",	
												x"074d",	x"0753",	x"072d",	x"0740",	
												x"0772",	x"072b",	x"0781",	x"0773",	
												x"0783",	x"075e",	x"0780",	x"0770",	
												x"0791",	x"0763",	x"07a0",	x"0765",	
												x"0779",	x"076d",	x"0718",	x"072a",	
												x"5031",	x"137c",	x"0728",	x"0706",	
												x"074f",	x"0726",	x"074d",	x"071b",	
												x"0742",	x"0707",	x"074c",	x"0722",	
												x"0752",	x"0713",	x"0745",	x"0718",	
												x"072b",	x"073b",	x"076f",	x"0721",	
												x"0789",	x"074a",	x"0780",	x"074e",	
												x"0775",	x"074e",	x"0774",	x"0770",	
												x"077a",	x"075c",	x"0773",	x"075b",	
												x"0768",	x"0756",	x"078c",	x"075b",	
												x"0792",	x"0774",	x"077d",	x"0765",	
												x"07aa",	x"076d",	x"07b0",	x"0747",	
												x"07a4",	x"0789",	x"07a2",	x"0772",	
												x"0784",	x"075a",	x"07ac",	x"0758",	
												x"07ba",	x"0798",	x"07c8",	x"0764",	
												x"07a9",	x"0792",	x"07b7",	x"0769",	
												x"07a9",	x"07a2",	x"079b",	x"077f",	
												x"0729",	x"076d",	x"6031",	x"137c",	
												x"074d",	x"0710",	x"075b",	x"073a",	
												x"074b",	x"0735",	x"0751",	x"0710",	
												x"0737",	x"0733",	x"0749",	x"0704",	
												x"0764",	x"06ff",	x"0742",	x"0725",	
												x"0795",	x"072e",	x"078d",	x"076b",	
												x"079a",	x"074a",	x"07cb",	x"0791",	
												x"07b6",	x"0792",	x"07b1",	x"078e",	
												x"07ce",	x"0775",	x"0794",	x"077a",	
												x"07bb",	x"078d",	x"07c6",	x"079b",	
												x"07cd",	x"079b",	x"07d3",	x"07bf",	
												x"07db",	x"07ae",	x"07e2",	x"07a6",	
												x"07b3",	x"07a9",	x"07ac",	x"079b",	
												x"07ee",	x"0788",	x"0803",	x"07c6",	
												x"07f5",	x"07ab",	x"0808",	x"07b9",	
												x"0801",	x"07c0",	x"0800",	x"07d4",	
												x"07e1",	x"07b6",	x"078b",	x"07a0",	
												x"7031",	x"137c",	x"07ac",	x"077b",	
												x"07c3",	x"0781",	x"07a5",	x"0799",	
												x"07c0",	x"079c",	x"07c5",	x"0774",	
												x"07a7",	x"0787",	x"079e",	x"0768",	
												x"07b0",	x"0799",	x"080b",	x"07a7",	
												x"0813",	x"07d6",	x"0822",	x"07c8",	
												x"081e",	x"0821",	x"0829",	x"0808",	
												x"085b",	x"0820",	x"0810",	x"080f",	
												x"081b",	x"0806",	x"0845",	x"07e7",	
												x"085f",	x"0816",	x"084e",	x"0816",	
												x"0841",	x"0822",	x"084b",	x"0825",	
												x"086a",	x"082e",	x"084e",	x"0846",	
												x"081a",	x"0835",	x"0869",	x"0833",	
												x"08b0",	x"0835",	x"088c",	x"0843",	
												x"087e",	x"0850",	x"08a5",	x"084f",	
												x"08a5",	x"0874",	x"0882",	x"0876",	
												x"076f",	x"084f",	x"0004",	x"000a",	
												x"6f64",	x"8f1c",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"237d",	
												x"0787",	x"079d",	x"0786",	x"0781",	
												x"071f",	x"0760",	x"0760",	x"0761",	
												x"075e",	x"075f",	x"0785",	x"075d",	
												x"0762",	x"0784",	x"078b",	x"0781",	
												x"078a",	x"0797",	x"0782",	x"078a",	
												x"079d",	x"0785",	x"0787",	x"078d",	
												x"0799",	x"0789",	x"0798",	x"077b",	
												x"07b3",	x"07bb",	x"0745",	x"078c",	
												x"0785",	x"0780",	x"0785",	x"0788",	
												x"079b",	x"076d",	x"0786",	x"0788",	
												x"07a9",	x"07ac",	x"07aa",	x"07aa",	
												x"07c9",	x"07c1",	x"079b",	x"07c2",	
												x"07a7",	x"077d",	x"07a3",	x"07a0",	
												x"07ba",	x"07b6",	x"0797",	x"07b7",	
												x"07a7",	x"078a",	x"07b6",	x"0792",	
												x"07bf",	x"078c",	x"0773",	x"07a7",	
												x"1031",	x"237d",	x"0759",	x"0778",	
												x"073d",	x"074f",	x"075e",	x"074b",	
												x"071c",	x"074d",	x"0754",	x"0750",	
												x"0796",	x"0739",	x"076b",	x"077c",	
												x"075f",	x"077d",	x"07af",	x"0768",	
												x"07a7",	x"079f",	x"07a0",	x"0787",	
												x"0771",	x"07be",	x"077b",	x"0789",	
												x"0794",	x"07a1",	x"0771",	x"07a1",	
												x"0770",	x"078d",	x"077c",	x"0795",	
												x"077e",	x"0784",	x"0771",	x"0779",	
												x"077a",	x"0793",	x"076c",	x"0788",	
												x"07a2",	x"0792",	x"0799",	x"0792",	
												x"0764",	x"07a3",	x"077c",	x"078c",	
												x"07c1",	x"07b7",	x"07a5",	x"07d1",	
												x"07ae",	x"0790",	x"07a9",	x"07c0",	
												x"07b2",	x"07b1",	x"07ae",	x"0796",	
												x"0745",	x"079b",	x"2031",	x"237d",	
												x"0759",	x"0759",	x"0728",	x"075e",	
												x"075e",	x"0738",	x"074c",	x"073e",	
												x"0749",	x"072b",	x"073c",	x"0747",	
												x"0776",	x"0762",	x"0712",	x"077d",	
												x"0779",	x"0746",	x"077c",	x"079a",	
												x"0769",	x"077c",	x"074e",	x"0763",	
												x"0782",	x"0769",	x"0780",	x"078d",	
												x"077c",	x"0772",	x"074d",	x"0769",	
												x"0761",	x"075a",	x"0790",	x"075c",	
												x"077f",	x"0788",	x"0762",	x"0776",	
												x"0779",	x"0766",	x"0780",	x"07a5",	
												x"0788",	x"077c",	x"077e",	x"076f",	
												x"07a5",	x"076a",	x"077d",	x"0770",	
												x"07a2",	x"077a",	x"077a",	x"0783",	
												x"078b",	x"0784",	x"0790",	x"0778",	
												x"0796",	x"0788",	x"071d",	x"076f",	
												x"3031",	x"237d",	x"0734",	x"072e",	
												x"074a",	x"0721",	x"0724",	x"0721",	
												x"0724",	x"071e",	x"071a",	x"06fe",	
												x"0741",	x"0725",	x"072f",	x"071e",	
												x"070f",	x"0720",	x"0777",	x"073b",	
												x"076e",	x"076d",	x"0764",	x"0764",	
												x"0766",	x"0754",	x"0773",	x"0743",	
												x"0777",	x"074f",	x"077d",	x"0772",	
												x"073f",	x"076f",	x"0766",	x"0763",	
												x"075a",	x"0784",	x"0768",	x"0756",	
												x"078a",	x"0761",	x"0794",	x"0768",	
												x"078f",	x"077f",	x"0793",	x"076c",	
												x"0772",	x"0777",	x"07bd",	x"074d",	
												x"0799",	x"077f",	x"0797",	x"077e",	
												x"0796",	x"0771",	x"07a9",	x"0777",	
												x"0798",	x"077b",	x"07aa",	x"0784",	
												x"073d",	x"0777",	x"0004",	x"000a",	
												x"5c0f",	x"cd43",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"237e",	
												x"0763",	x"0754",	x"074f",	x"0714",	
												x"0753",	x"073b",	x"0741",	x"0754",	
												x"075b",	x"073f",	x"076c",	x"076d",	
												x"0764",	x"0757",	x"0763",	x"0757",	
												x"079c",	x"076d",	x"078a",	x"077b",	
												x"078a",	x"077e",	x"0793",	x"077e",	
												x"0792",	x"0781",	x"07d0",	x"0798",	
												x"07a3",	x"0798",	x"079e",	x"0787",	
												x"07af",	x"07ac",	x"07a9",	x"07ae",	
												x"07d1",	x"07ca",	x"07be",	x"07b0",	
												x"07c1",	x"07ba",	x"07c8",	x"07b0",	
												x"07e7",	x"07c4",	x"07c0",	x"07d7",	
												x"07eb",	x"07c8",	x"07d5",	x"07c5",	
												x"07d8",	x"07cb",	x"07c8",	x"07df",	
												x"07eb",	x"07cc",	x"07d3",	x"07d0",	
												x"07db",	x"07c4",	x"077c",	x"07df",	
												x"5031",	x"237e",	x"0791",	x"0778",	
												x"0798",	x"0789",	x"0797",	x"075d",	
												x"07c6",	x"0790",	x"07b7",	x"077b",	
												x"07ba",	x"077f",	x"07ce",	x"07a1",	
												x"07a1",	x"079a",	x"07e5",	x"0791",	
												x"07f3",	x"07cc",	x"07e4",	x"07cd",	
												x"080b",	x"07d3",	x"07ef",	x"07cf",	
												x"080d",	x"07da",	x"07f9",	x"07dc",	
												x"07f5",	x"07d2",	x"07ef",	x"07a8",	
												x"080e",	x"07b1",	x"080e",	x"07b6",	
												x"0822",	x"07ef",	x"081c",	x"07e7",	
												x"0827",	x"07f3",	x"0827",	x"07fe",	
												x"07fd",	x"0809",	x"0839",	x"07e3",	
												x"082f",	x"07da",	x"082a",	x"07e7",	
												x"0831",	x"07f1",	x"083f",	x"07e5",	
												x"0835",	x"0813",	x"0821",	x"080b",	
												x"0795",	x"07e4",	x"6031",	x"237e",	
												x"07a3",	x"0783",	x"079f",	x"0788",	
												x"07bb",	x"0776",	x"07e3",	x"077d",	
												x"07b1",	x"0793",	x"07d5",	x"077f",	
												x"07d6",	x"07ba",	x"07cd",	x"07b5",	
												x"07fc",	x"07c7",	x"0818",	x"07f4",	
												x"0825",	x"07d7",	x"084e",	x"07e8",	
												x"083d",	x"07e6",	x"0822",	x"07ea",	
												x"083d",	x"07f9",	x"0837",	x"07e7",	
												x"0820",	x"07f9",	x"0841",	x"0810",	
												x"084f",	x"0811",	x"0853",	x"081d",	
												x"0897",	x"0821",	x"088e",	x"0829",	
												x"0851",	x"0837",	x"0861",	x"082a",	
												x"085d",	x"0832",	x"0842",	x"0838",	
												x"085f",	x"082f",	x"086a",	x"0823",	
												x"0868",	x"080c",	x"086f",	x"0834",	
												x"0857",	x"082d",	x"07fc",	x"0838",	
												x"7031",	x"237e",	x"0819",	x"07d9",	
												x"0825",	x"0809",	x"0842",	x"07cb",	
												x"0840",	x"07d1",	x"082c",	x"07f7",	
												x"0862",	x"0812",	x"0883",	x"081c",	
												x"0841",	x"082f",	x"0882",	x"083c",	
												x"089b",	x"086f",	x"0898",	x"088e",	
												x"08a4",	x"086a",	x"089f",	x"0868",	
												x"08b1",	x"0880",	x"08ad",	x"0894",	
												x"0888",	x"0877",	x"08ba",	x"086a",	
												x"08ce",	x"089e",	x"08c0",	x"0892",	
												x"08d1",	x"0893",	x"08d2",	x"0895",	
												x"08d6",	x"08c7",	x"08ce",	x"08cc",	
												x"08c8",	x"08d3",	x"08e4",	x"08c4",	
												x"08d6",	x"08ca",	x"08ea",	x"08bc",	
												x"08fb",	x"08cf",	x"0906",	x"08a6",	
												x"0910",	x"08db",	x"08f3",	x"08df",	
												x"0702",	x"08e5",	x"0004",	x"000a",	
												x"aa3e",	x"0a50",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"0031",	x"337f",	
												x"06b0",	x"0713",	x"06cd",	x"06a0",	
												x"06a3",	x"06b7",	x"06b6",	x"068a",	
												x"06ac",	x"06be",	x"06c8",	x"06c5",	
												x"06ac",	x"06c3",	x"06a8",	x"06b8",	
												x"06f3",	x"06b4",	x"06e7",	x"0701",	
												x"06e3",	x"071a",	x"0700",	x"071a",	
												x"06ea",	x"06f7",	x"0701",	x"0720",	
												x"06ef",	x"0715",	x"06bf",	x"06ea",	
												x"06ec",	x"06fb",	x"070a",	x"06f2",	
												x"0703",	x"0716",	x"06e9",	x"0705",	
												x"06f5",	x"0700",	x"0700",	x"06fb",	
												x"06f1",	x"0712",	x"06dc",	x"0734",	
												x"06eb",	x"0702",	x"070b",	x"0705",	
												x"070e",	x"0710",	x"06e4",	x"0708",	
												x"06e6",	x"070f",	x"072a",	x"06f2",	
												x"070d",	x"0710",	x"06b9",	x"0704",	
												x"1031",	x"337f",	x"06ce",	x"06a5",	
												x"06b1",	x"06bf",	x"069f",	x"06a7",	
												x"06a6",	x"06a0",	x"06a2",	x"06a1",	
												x"0699",	x"06af",	x"06eb",	x"06c8",	
												x"069c",	x"06e4",	x"06cb",	x"06b9",	
												x"06f0",	x"06e5",	x"06e9",	x"06e0",	
												x"06dc",	x"06dc",	x"06db",	x"06d2",	
												x"06f0",	x"06f0",	x"06c3",	x"06df",	
												x"06c0",	x"06be",	x"06f0",	x"06db",	
												x"06d7",	x"070a",	x"06d9",	x"06f4",	
												x"06e5",	x"06fd",	x"06da",	x"06fd",	
												x"071b",	x"06fc",	x"0717",	x"0704",	
												x"06ca",	x"070b",	x"06fd",	x"06d8",	
												x"0704",	x"0708",	x"06ef",	x"06fa",	
												x"0710",	x"070d",	x"06fb",	x"0708",	
												x"072c",	x"06f7",	x"0719",	x"070d",	
												x"06bd",	x"0709",	x"2031",	x"337f",	
												x"06c5",	x"06bc",	x"06aa",	x"06cf",	
												x"06c7",	x"06a5",	x"0690",	x"06ae",	
												x"069c",	x"0694",	x"06af",	x"06a3",	
												x"06b5",	x"06c7",	x"06ad",	x"06dd",	
												x"06db",	x"06c3",	x"06db",	x"06e6",	
												x"06dd",	x"06ec",	x"06c8",	x"06fa",	
												x"06dd",	x"06de",	x"06e8",	x"06ef",	
												x"06f0",	x"06e6",	x"06b5",	x"06e3",	
												x"06ea",	x"06c3",	x"0703",	x"06e1",	
												x"06e0",	x"06e8",	x"06da",	x"06d8",	
												x"06d2",	x"06d5",	x"06e9",	x"06d0",	
												x"06d8",	x"06f0",	x"06d0",	x"06c7",	
												x"070c",	x"06e5",	x"06f0",	x"0700",	
												x"06f0",	x"06e7",	x"06f2",	x"06be",	
												x"06ef",	x"06d5",	x"06fb",	x"06e7",	
												x"06fa",	x"06db",	x"06bb",	x"06e3",	
												x"3031",	x"337f",	x"068f",	x"06b2",	
												x"068c",	x"0693",	x"06a8",	x"066b",	
												x"06bf",	x"067f",	x"0676",	x"066f",	
												x"06c0",	x"0680",	x"069d",	x"06b0",	
												x"06a2",	x"068c",	x"06ba",	x"06ae",	
												x"06d7",	x"06b5",	x"06e0",	x"06a8",	
												x"06e0",	x"06d0",	x"06dc",	x"06d1",	
												x"06d5",	x"06c3",	x"06dc",	x"06c7",	
												x"06cc",	x"06d5",	x"06db",	x"06ac",	
												x"06e7",	x"06d0",	x"06f8",	x"06dd",	
												x"06fd",	x"06eb",	x"06e6",	x"06e3",	
												x"0714",	x"06f5",	x"0709",	x"06ef",	
												x"06f5",	x"06d1",	x"0701",	x"06d8",	
												x"06fc",	x"06e7",	x"06ff",	x"06dd",	
												x"070d",	x"06ee",	x"071c",	x"06eb",	
												x"0709",	x"06cb",	x"070c",	x"06ee",	
												x"06b4",	x"06e5",	x"0004",	x"000a",	
												x"0d9f",	x"bf89",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"ffee",	x"00c0",	
												x"d125",	x"0000",	x"4031",	x"3380",	
												x"06b9",	x"06a0",	x"06cd",	x"067a",	
												x"06d5",	x"0681",	x"06db",	x"069e",	
												x"06cd",	x"0699",	x"06f4",	x"06a8",	
												x"06c3",	x"06ba",	x"06cf",	x"06a7",	
												x"0704",	x"06cf",	x"0712",	x"06e8",	
												x"06ff",	x"0702",	x"06f7",	x"06fb",	
												x"071c",	x"06e6",	x"070f",	x"0703",	
												x"0710",	x"070a",	x"06f5",	x"0715",	
												x"0732",	x"06f8",	x"0709",	x"071b",	
												x"0725",	x"0708",	x"0726",	x"0732",	
												x"0735",	x"0728",	x"073c",	x"071b",	
												x"074c",	x"0710",	x"0735",	x"0728",	
												x"0732",	x"071c",	x"0731",	x"0714",	
												x"073e",	x"071b",	x"073e",	x"071d",	
												x"075b",	x"072c",	x"077a",	x"0745",	
												x"074a",	x"0740",	x"06e8",	x"071d",	
												x"5031",	x"3380",	x"072e",	x"06f6",	
												x"06fc",	x"06dd",	x"06fc",	x"06b3",	
												x"06f9",	x"06c9",	x"06f5",	x"06d8",	
												x"0722",	x"06d2",	x"0712",	x"0710",	
												x"0709",	x"06ee",	x"0739",	x"0701",	
												x"073d",	x"0720",	x"0744",	x"0736",	
												x"073b",	x"0739",	x"075d",	x"0730",	
												x"0742",	x"0745",	x"0742",	x"0728",	
												x"0727",	x"0740",	x"074a",	x"0720",	
												x"0756",	x"0739",	x"075d",	x"073a",	
												x"0774",	x"0758",	x"079b",	x"0750",	
												x"0784",	x"0740",	x"0779",	x"0743",	
												x"0762",	x"0740",	x"0799",	x"0743",	
												x"0784",	x"0750",	x"077d",	x"074d",	
												x"076e",	x"074b",	x"0782",	x"0741",	
												x"07c5",	x"0756",	x"0777",	x"074e",	
												x"0709",	x"0762",	x"6031",	x"3380",	
												x"071d",	x"06fd",	x"0717",	x"06f4",	
												x"070a",	x"06e3",	x"0719",	x"06de",	
												x"0711",	x"06f4",	x"073d",	x"070d",	
												x"073c",	x"0712",	x"073f",	x"0741",	
												x"075f",	x"072c",	x"0790",	x"073f",	
												x"0777",	x"075b",	x"077b",	x"0754",	
												x"076e",	x"0769",	x"079c",	x"0772",	
												x"0798",	x"0770",	x"0779",	x"075f",	
												x"0779",	x"0757",	x"078b",	x"0783",	
												x"0794",	x"077b",	x"07b4",	x"078f",	
												x"0789",	x"076a",	x"07a2",	x"077e",	
												x"07c8",	x"0780",	x"07a2",	x"0790",	
												x"07d4",	x"076e",	x"07c8",	x"079a",	
												x"07d0",	x"078a",	x"07d7",	x"0797",	
												x"07dc",	x"078f",	x"07d8",	x"07ac",	
												x"07b3",	x"07a4",	x"074c",	x"077f",	
												x"7031",	x"3380",	x"0773",	x"0754",	
												x"079a",	x"075b",	x"0767",	x"0734",	
												x"07bf",	x"071e",	x"079f",	x"0724",	
												x"07a4",	x"0761",	x"0791",	x"0763",	
												x"078c",	x"0768",	x"07ee",	x"076d",	
												x"07f6",	x"07af",	x"07e2",	x"07c2",	
												x"07fa",	x"07ba",	x"07ec",	x"07a7",	
												x"07f3",	x"07d4",	x"07f2",	x"07b1",	
												x"07f2",	x"07cc",	x"080f",	x"07cb",	
												x"081f",	x"07f8",	x"07fd",	x"07cf",	
												x"0808",	x"07f7",	x"0811",	x"0800",	
												x"0823",	x"07fd",	x"081a",	x"07fc",	
												x"0808",	x"07f6",	x"083e",	x"0802",	
												x"0816",	x"081a",	x"0865",	x"07f3",	
												x"0856",	x"0818",	x"085e",	x"0806",	
												x"085e",	x"0820",	x"084c",	x"082e",	
												x"0742",	x"0814",	x"0004",	x"000a",	
												x"5936",	x"f86e",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"b10c",	x"ce11",	
												x"d125",	x"0000",	x"0000",	x"0081",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"0004",	x"000a",	
												x"bcc5",	x"1e89",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"b0de",	x"000a",	
												x"d125",	x"0000",	x"0000",	x"0082",	
												x"03e8",	x"03e8",	x"03e8",	x"03e8",	
												x"03e8",	x"03e8",	x"03e8",	x"03e8",	
												x"03e8",	x"03e8",	x"03e8",	x"03e8",	
												x"03e8",	x"03e8",	x"03e8",	x"03e8",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"079e",	x"079e",	x"079e",	x"079e",	
												x"051e",	x"051e",	x"051e",	x"051e",	
												x"051e",	x"051e",	x"051e",	x"051e",	
												x"051e",	x"051e",	x"051e",	x"051e",	
												x"051e",	x"051e",	x"051e",	x"051e",	
												x"0c9e",	x"0c9e",	x"0c9e",	x"0c9e",	
												x"0c9e",	x"0c9e",	x"0c9e",	x"0c9e",	
												x"0c9e",	x"0c9e",	x"0c9e",	x"0c9e",	
												x"0c9e",	x"0c9e",	x"0c9e",	x"0c9e",	
												x"042e",	x"042e",	x"042e",	x"042e",	
												x"042e",	x"042e",	x"042e",	x"042e",	
												x"042e",	x"042e",	x"042e",	x"042e",	
												x"042e",	x"042e",	x"042e",	x"042e",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"0640",	x"0640",	x"0640",	x"0640",	
												x"0640",	x"0640",	x"0640",	x"0640",	
												x"0640",	x"0640",	x"0640",	x"0640",	
												x"0640",	x"0640",	x"0640",	x"0640",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"044c",	x"044c",	x"044c",	x"044c",	
												x"0883",	x"0913",	x"09c8",	x"09a9",	
												x"085a",	x"09ea",	x"099d",	x"08de",	
												x"0e7a",	x"0a2f",	x"0c8b",	x"0c45",	
												x"0afd",	x"0c7c",	x"0e24",	x"0982",	
												x"0384",	x"0384",	x"0384",	x"0384",	
												x"0384",	x"0384",	x"0384",	x"0384",	
												x"0384",	x"0384",	x"0384",	x"0384",	
												x"0384",	x"0384",	x"0384",	x"0384",	
												x"0ce4",	x"0ce4",	x"0ce4",	x"0ce4",	
												x"0ce4",	x"0ce4",	x"0ce4",	x"0ce4",	
												x"0ce4",	x"0ce4",	x"0ce4",	x"0ce4",	
												x"0ce4",	x"0ce4",	x"0ce4",	x"0ce4",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"050f",	x"0000",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"0004",	x"000a",	
												x"098d",	x"9200",	x"4944",	x"6250",	
												x"11e2",	x"00be",	x"008c",	x"0000",	
												x"1213",	x"2011",	x"00da",	x"000f",	
												x"d125",	x"0000",	x"0000",	x"0083",	
												x"ffff",	x"0000",	x"079d",	x"0000",	
												x"079c",	x"0000",	x"079e",	x"0000",	
												x"079d",	x"0000",	x"07a8",	x"0000",	
												x"079c",	x"0000",	x"079e",	x"0000",	
												x"07a1",	x"0000",	x"079d",	x"0000",	
												x"079c",	x"0000",	x"079c",	x"0000",	
												x"079c",	x"0000",	x"079d",	x"0000",	
												x"079d",	x"0000",	x"079d",	x"0000",	
												x"0799",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"0000",	x"0000",	x"0000",	x"0000",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"9999",	x"9999",	
												x"9999",	x"9999",	x"0004",	x"000a",	
												x"ec98",	x"b6f0",	x"4944",	x"6250"
										);
end data16_pkg;